// Tom has a total of 208 pins, taken from the schematic by Atari:
// 14 input  pins VCC
// 24 input  pins GND
// 64 inout  pins data bus
// 24 inout  pins address bus
// 11 inout  pins are MA
// 3  inout  pins are FC
// 2  inout  pins are SIZ
// 8  output pins Red
// 8  output pins Green
// 8  output pins Blue
// 2  output Pins DBRL
// 2  output Pins ROMCSL
// 2  output pins RAS
// 2  output pins CAS
// 2  output pins OEL
// 8  output pins WEL
// 3  output pins MASKA
// 1  output pin HSL (Hsync)
// 1  output pin VSL (Vsync)
// 1  output pin LP
// 1  output pin Inc
// 1  output pin DREOL
// 1  output pin DTACKL
// 1  output pin RW
// 1  output pin INTL
// 1  output pin DINT
// 1  output pin BRL
// 1  output pin BGL
// 1  output pin BGA
// 1  output pin DSPCSL
// 1  output pin RESETL
// 1  output pin TEST
// 1  output pin VCLK -- "20 mil trooo(?) on clocks" -- pclkosc on jerry, 26.6mhz
// 1  output pin PCLK -- sysclk on jerry
// 1  output pin WAITL
// 1  output pin EXPL

module tom_w (
	// Real Pins. Inout pins have been split.
	output [63:0]  dbus_out,
	input  [63:0]  dbus_in,
	output [23:0]  abus_out,
	input  [23:0]  abus_in,
	output [10:0]  MA_out,
	input  [10:0]  MA_in,
	output [2:0]   FC_out,
	input  [2:0]   FC_in,
	output [1:0]   SIZ_out,
	input  [1:0]   SIZ_in,
	output [8:0]   red,
	output [8:0]   green,
	output [8:0]   blue,
	input  [1:0]   DBR_n,
	output [1:0]   ROM_CS_n,
	output [1:0]   RAS,
	output [1:0]   CAS,
	output [1:0]   OE_n,
	output [7:0]   WE_n,
	output [2:0]   MASKA,
	output         HS_out_n,
	input          HS_in_n,
	output         VS_out_n,
	input          VS_in_n,
	input          LP,
	output         INC,
	output         DREO_n,
	output         DTACK_n,
	output         RW,
	output         INT_n,
	input          DINT,
	output         BR_n,
	output         BG_n,
	output         BGA_out, // BA?
	input          BGA_in, // BA?
	output         DSP_CS_n,
	input          RESET_n,
	input          TEST,
	input          VCLK,
	input          PCLK,
	input          WAIT_n,
	output         EXP_n,
	// Abstracted Pins to assist with FPGA implementation
	output [63:0]  dbus_oe, // Indicates that a particular data pins output is driven
	input  [23:0]  abus_oe,
	output [10:0]  MA_oe,
	output [1:0]   SIZ_oe,
	output         BGA_oe, // BA?
	output [1:0]   DBR_oe,
	output         HS_oe,
	// Completely 
	input          clk_sys,
	input          ram_ready,
	input          tlw // This appears to be a signal to indicate the address bus is ready to latch
);

// TOM
tom tom_inst
(
	.xbgl(xbgl),
	.xdbrl_0(xdbrl[0]),
	.xdbrl_1(xdbrl[1]),
	.xlp(xlp),
	.xdint(xdint),
	.xtest(xtest),
	.xpclk(xpclk),
	.xvclk(xvclk),
	.xwaitl(xwaitl),
	.xresetl(xresetl),
	.xd_0_out(dbus_out[0]),
	.xd_0_oe(dbus_oe[0]),
	.xd_0_in(dbus_in[0]),
	.xd_1_out(dbus_out[1]),
	.xd_1_oe(dbus_oe[1]),
	.xd_1_in(dbus_in[1]),
	.xd_2_out(dbus_out[2]),
	.xd_2_oe(dbus_oe[2]),
	.xd_2_in(dbus_in[2]),
	.xd_3_out(dbus_out[3]),
	.xd_3_oe(dbus_oe[3]),
	.xd_3_in(dbus_in[3]),
	.xd_4_out(dbus_out[4]),
	.xd_4_oe(dbus_oe[4]),
	.xd_4_in(dbus_in[4]),
	.xd_5_out(dbus_out[5]),
	.xd_5_oe(dbus_oe[5]),
	.xd_5_in(dbus_in[5]),
	.xd_6_out(dbus_out[6]),
	.xd_6_oe(dbus_oe[6]),
	.xd_6_in(dbus_in[6]),
	.xd_7_out(dbus_out[7]),
	.xd_7_oe(dbus_oe[7]),
	.xd_7_in(dbus_in[7]),
	.xd_8_out(dbus_out[8]),
	.xd_8_oe(dbus_oe[8]),
	.xd_8_in(dbus_in[8]),
	.xd_9_out(dbus_out[9]),
	.xd_9_oe(dbus_oe[9]),
	.xd_9_in(dbus_in[9]),
	.xd_10_out(dbus_out[10]),
	.xd_10_oe(dbus_oe[10]),
	.xd_10_in(dbus_in[10]),
	.xd_11_out(dbus_out[11]),
	.xd_11_oe(dbus_oe[11]),
	.xd_11_in(dbus_in[11]),
	.xd_12_out(dbus_out[12]),
	.xd_12_oe(dbus_oe[12]),
	.xd_12_in(dbus_in[12]),
	.xd_13_out(dbus_out[13]),
	.xd_13_oe(dbus_oe[13]),
	.xd_13_in(dbus_in[13]),
	.xd_14_out(dbus_out[14]),
	.xd_14_oe(dbus_oe[14]),
	.xd_14_in(dbus_in[14]),
	.xd_15_out(dbus_out[15]),
	.xd_15_oe(dbus_oe[15]),
	.xd_15_in(dbus_in[15]),
	.xd_16_out(dbus_out[16]),
	.xd_16_oe(dbus_oe[16]),
	.xd_16_in(dbus_in[16]),
	.xd_17_out(dbus_out[17]),
	.xd_17_oe(dbus_oe[17]),
	.xd_17_in(dbus_in[17]),
	.xd_18_out(dbus_out[18]),
	.xd_18_oe(dbus_oe[18]),
	.xd_18_in(dbus_in[18]),
	.xd_19_out(dbus_out[19]),
	.xd_19_oe(dbus_oe[19]),
	.xd_19_in(dbus_in[19]),
	.xd_20_out(dbus_out[20]),
	.xd_20_oe(dbus_oe[20]),
	.xd_20_in(dbus_in[20]),
	.xd_21_out(dbus_out[21]),
	.xd_21_oe(dbus_oe[21]),
	.xd_21_in(dbus_in[21]),
	.xd_22_out(dbus_out[22]),
	.xd_22_oe(dbus_oe[22]),
	.xd_22_in(dbus_in[22]),
	.xd_23_out(dbus_out[23]),
	.xd_23_oe(dbus_oe[23]),
	.xd_23_in(dbus_in[23]),
	.xd_24_out(dbus_out[24]),
	.xd_24_oe(dbus_oe[24]),
	.xd_24_in(dbus_in[24]),
	.xd_25_out(dbus_out[25]),
	.xd_25_oe(dbus_oe[25]),
	.xd_25_in(dbus_in[25]),
	.xd_26_out(dbus_out[26]),
	.xd_26_oe(dbus_oe[26]),
	.xd_26_in(dbus_in[26]),
	.xd_27_out(dbus_out[27]),
	.xd_27_oe(dbus_oe[27]),
	.xd_27_in(dbus_in[27]),
	.xd_28_out(dbus_out[28]),
	.xd_28_oe(dbus_oe[28]),
	.xd_28_in(dbus_in[28]),
	.xd_29_out(dbus_out[29]),
	.xd_29_oe(dbus_oe[29]),
	.xd_29_in(dbus_in[29]),
	.xd_30_out(dbus_out[30]),
	.xd_30_oe(dbus_oe[30]),
	.xd_30_in(dbus_in[30]),
	.xd_31_out(dbus_out[31]),
	.xd_31_oe(dbus_oe[31]),
	.xd_31_in(dbus_in[31]),
	.xd_32_out(dbus_out[32]),
	.xd_32_oe(dbus_oe[32]),
	.xd_32_in(dbus_in[32]),
	.xd_33_out(dbus_out[33]),
	.xd_33_oe(dbus_oe[33]),
	.xd_33_in(dbus_in[33]),
	.xd_34_out(dbus_out[34]),
	.xd_34_oe(dbus_oe[34]),
	.xd_34_in(dbus_in[34]),
	.xd_35_out(dbus_out[35]),
	.xd_35_oe(dbus_oe[35]),
	.xd_35_in(dbus_in[35]),
	.xd_36_out(dbus_out[36]),
	.xd_36_oe(dbus_oe[36]),
	.xd_36_in(dbus_in[36]),
	.xd_37_out(dbus_out[37]),
	.xd_37_oe(dbus_oe[37]),
	.xd_37_in(dbus_in[37]),
	.xd_38_out(dbus_out[38]),
	.xd_38_oe(dbus_oe[38]),
	.xd_38_in(dbus_in[38]),
	.xd_39_out(dbus_out[39]),
	.xd_39_oe(dbus_oe[39]),
	.xd_39_in(dbus_in[39]),
	.xd_40_out(dbus_out[40]),
	.xd_40_oe(dbus_oe[40]),
	.xd_40_in(dbus_in[40]),
	.xd_41_out(dbus_out[41]),
	.xd_41_oe(dbus_oe[41]),
	.xd_41_in(dbus_in[41]),
	.xd_42_out(dbus_out[42]),
	.xd_42_oe(dbus_oe[42]),
	.xd_42_in(dbus_in[42]),
	.xd_43_out(dbus_out[43]),
	.xd_43_oe(dbus_oe[43]),
	.xd_43_in(dbus_in[43]),
	.xd_44_out(dbus_out[44]),
	.xd_44_oe(dbus_oe[44]),
	.xd_44_in(dbus_in[44]),
	.xd_45_out(dbus_out[45]),
	.xd_45_oe(dbus_oe[45]),
	.xd_45_in(dbus_in[45]),
	.xd_46_out(dbus_out[46]),
	.xd_46_oe(dbus_oe[46]),
	.xd_46_in(dbus_in[46]),
	.xd_47_out(dbus_out[47]),
	.xd_47_oe(dbus_oe[47]),
	.xd_47_in(dbus_in[47]),
	.xd_48_out(dbus_out[48]),
	.xd_48_oe(dbus_oe[48]),
	.xd_48_in(dbus_in[48]),
	.xd_49_out(dbus_out[49]),
	.xd_49_oe(dbus_oe[49]),
	.xd_49_in(dbus_in[49]),
	.xd_50_out(dbus_out[50]),
	.xd_50_oe(dbus_oe[50]),
	.xd_50_in(dbus_in[50]),
	.xd_51_out(dbus_out[51]),
	.xd_51_oe(dbus_oe[51]),
	.xd_51_in(dbus_in[51]),
	.xd_52_out(dbus_out[52]),
	.xd_52_oe(dbus_oe[52]),
	.xd_52_in(dbus_in[52]),
	.xd_53_out(dbus_out[53]),
	.xd_53_oe(dbus_oe[53]),
	.xd_53_in(dbus_in[53]),
	.xd_54_out(dbus_out[54]),
	.xd_54_oe(dbus_oe[54]),
	.xd_54_in(dbus_in[54]),
	.xd_55_out(dbus_out[55]),
	.xd_55_oe(dbus_oe[55]),
	.xd_55_in(dbus_in[55]),
	.xd_56_out(dbus_out[56]),
	.xd_56_oe(dbus_oe[56]),
	.xd_56_in(dbus_in[56]),
	.xd_57_out(dbus_out[57]),
	.xd_57_oe(dbus_oe[57]),
	.xd_57_in(dbus_in[57]),
	.xd_58_out(dbus_out[58]),
	.xd_58_oe(dbus_oe[58]),
	.xd_58_in(dbus_in[58]),
	.xd_59_out(dbus_out[59]),
	.xd_59_oe(dbus_oe[59]),
	.xd_59_in(dbus_in[59]),
	.xd_60_out(dbus_out[60]),
	.xd_60_oe(dbus_oe[60]),
	.xd_60_in(dbus_in[60]),
	.xd_61_out(dbus_out[61]),
	.xd_61_oe(dbus_oe[61]),
	.xd_61_in(dbus_in[61]),
	.xd_62_out(dbus_out[62]),
	.xd_62_oe(dbus_oe[62]),
	.xd_62_in(dbus_in[62]),
	.xd_63_out(dbus_out[63]),
	.xd_63_oe(dbus_oe[63]),
	.xd_63_in(dbus_in[63]),
	.xa_0_out(xa_out[0]),
	.xa_0_oe(xa_oe[0]),
	.xa_0_in(xa_in[0]),
	.xa_1_out(xa_out[1]),
	.xa_1_oe(xa_oe[1]),
	.xa_1_in(xa_in[1]),
	.xa_2_out(xa_out[2]),
	.xa_2_oe(xa_oe[2]),
	.xa_2_in(xa_in[2]),
	.xa_3_out(xa_out[3]),
	.xa_3_oe(xa_oe[3]),
	.xa_3_in(xa_in[3]),
	.xa_4_out(xa_out[4]),
	.xa_4_oe(xa_oe[4]),
	.xa_4_in(xa_in[4]),
	.xa_5_out(xa_out[5]),
	.xa_5_oe(xa_oe[5]),
	.xa_5_in(xa_in[5]),
	.xa_6_out(xa_out[6]),
	.xa_6_oe(xa_oe[6]),
	.xa_6_in(xa_in[6]),
	.xa_7_out(xa_out[7]),
	.xa_7_oe(xa_oe[7]),
	.xa_7_in(xa_in[7]),
	.xa_8_out(xa_out[8]),
	.xa_8_oe(xa_oe[8]),
	.xa_8_in(xa_in[8]),
	.xa_9_out(xa_out[9]),
	.xa_9_oe(xa_oe[9]),
	.xa_9_in(xa_in[9]),
	.xa_10_out(xa_out[10]),
	.xa_10_oe(xa_oe[10]),
	.xa_10_in(xa_in[10]),
	.xa_11_out(xa_out[11]),
	.xa_11_oe(xa_oe[11]),
	.xa_11_in(xa_in[11]),
	.xa_12_out(xa_out[12]),
	.xa_12_oe(xa_oe[12]),
	.xa_12_in(xa_in[12]),
	.xa_13_out(xa_out[13]),
	.xa_13_oe(xa_oe[13]),
	.xa_13_in(xa_in[13]),
	.xa_14_out(xa_out[14]),
	.xa_14_oe(xa_oe[14]),
	.xa_14_in(xa_in[14]),
	.xa_15_out(xa_out[15]),
	.xa_15_oe(xa_oe[15]),
	.xa_15_in(xa_in[15]),
	.xa_16_out(xa_out[16]),
	.xa_16_oe(xa_oe[16]),
	.xa_16_in(xa_in[16]),
	.xa_17_out(xa_out[17]),
	.xa_17_oe(xa_oe[17]),
	.xa_17_in(xa_in[17]),
	.xa_18_out(xa_out[18]),
	.xa_18_oe(xa_oe[18]),
	.xa_18_in(xa_in[18]),
	.xa_19_out(xa_out[19]),
	.xa_19_oe(xa_oe[19]),
	.xa_19_in(xa_in[19]),
	.xa_20_out(xa_out[20]),
	.xa_20_oe(xa_oe[20]),
	.xa_20_in(xa_in[20]),
	.xa_21_out(xa_out[21]),
	.xa_21_oe(xa_oe[21]),
	.xa_21_in(xa_in[21]),
	.xa_22_out(xa_out[22]),
	.xa_22_oe(xa_oe[22]),
	.xa_22_in(xa_in[22]),
	.xa_23_out(xa_out[23]),
	.xa_23_oe(xa_oe[23]),
	.xa_23_in(xa_in[23]),
	.xma_0_out(xma_out[0]),
	.xma_0_oe(xma_oe[0]),
	.xma_0_in(xma_in[0]),
	.xma_1_out(xma_out[1]),
	.xma_1_oe(xma_oe[1]),
	.xma_1_in(xma_in[1]),
	.xma_2_out(xma_out[2]),
	.xma_2_oe(xma_oe[2]),
	.xma_2_in(xma_in[2]),
	.xma_3_out(xma_out[3]),
	.xma_3_oe(xma_oe[3]),
	.xma_3_in(xma_in[3]),
	.xma_4_out(xma_out[4]),
	.xma_4_oe(xma_oe[4]),
	.xma_4_in(xma_in[4]),
	.xma_5_out(xma_out[5]),
	.xma_5_oe(xma_oe[5]),
	.xma_5_in(xma_in[5]),
	.xma_6_out(xma_out[6]),
	.xma_6_oe(xma_oe[6]),
	.xma_6_in(xma_in[6]),
	.xma_7_out(xma_out[7]),
	.xma_7_oe(xma_oe[7]),
	.xma_7_in(xma_in[7]),
	.xma_8_out(xma_out[8]),
	.xma_8_oe(xma_oe[8]),
	.xma_8_in(xma_in[8]),
	.xma_9_out(xma_out[9]),
	.xma_9_oe(xma_oe[9]),
	.xma_9_in(xma_in[9]),
	.xma_10_out(xma_out[10]),
	.xma_10_oe(xma_oe[10]),
	.xma_10_in(xma_in[10]),
	.xhs_out(xhs_out),
	.xhs_oe(xhs_oe),
	.xhs_in(xhs_in),
	.xvs_out(xvs_out),
	.xvs_oe(xvs_oe),
	.xvs_in(xvs_in),
	.xsiz_0_out(xsiz_out[0]),
	.xsiz_0_oe(xsiz_oe[0]),
	.xsiz_0_in(xsiz_in[0]),
	.xsiz_1_out(xsiz_out[1]),
	.xsiz_1_oe(xsiz_oe[1]),
	.xsiz_1_in(xsiz_in[1]),
	.xfc_0_out(xfc_out[0]),
	.xfc_0_oe(xfc_oe[0]),
	.xfc_0_in(xfc_in[0]),
	.xfc_1_out(xfc_out[1]),
	.xfc_1_oe(xfc_oe[1]),
	.xfc_1_in(xfc_in[1]),
	.xfc_2_out(xfc_out[2]),
	.xfc_2_oe(xfc_oe[2]),
	.xfc_2_in(xfc_in[2]),
	.xrw_out(xrw_out),
	.xrw_oe(xrw_oe),
	.xrw_in(xrw_in),
	.xdreql_out(xdreql_out),
	.xdreql_oe(xdreql_oe),
	.xdreql_in(xdreql_in),
	.xba_out(xba_out),
	.xba_oe(xba_oe),
	.xba_in(xba_in),
	.xbrl_out(xbrl_out),
	.xbrl_oe(xbrl_oe),
	.xbrl_in(xbrl_in),
	.xr_0(xr[0]),
	.xr_1(xr[1]),
	.xr_2(xr[2]),
	.xr_3(xr[3]),
	.xr_4(xr[4]),
	.xr_5(xr[5]),
	.xr_6(xr[6]),
	.xr_7(xr[7]),
	.xg_0(xg[0]),
	.xg_1(xg[1]),
	.xg_2(xg[2]),
	.xg_3(xg[3]),
	.xg_4(xg[4]),
	.xg_5(xg[5]),
	.xg_6(xg[6]),
	.xg_7(xg[7]),
	.xb_0(xb[0]),
	.xb_1(xb[1]),
	.xb_2(xb[2]),
	.xb_3(xb[3]),
	.xb_4(xb[4]),
	.xb_5(xb[5]),
	.xb_6(xb[6]),
	.xb_7(xb[7]),
	.xinc(xinc),
	.xoel_0(xoel[0]),
	.xoel_1(xoel[1]),
	.xoel_2(xoel[2]),
	.xmaska_0(xmaska[0]),
	.xmaska_1(xmaska[1]),
	.xmaska_2(xmaska[2]),
	.xromcsl_0(xromcsl[0]),
	.xromcsl_1(xromcsl[1]),
	.xcasl_0(xcasl[0]),
	.xcasl_1(xcasl[1]),
	.xdbgl(xdbgl),
	.xexpl(xexpl),
	.xdspcsl(xdspcsl),
	.xwel_0(xwel[0]),
	.xwel_1(xwel[1]),
	.xwel_2(xwel[2]),
	.xwel_3(xwel[3]),
	.xwel_4(xwel[4]),
	.xwel_5(xwel[5]),
	.xwel_6(xwel[6]),
	.xwel_7(xwel[7]),
	.xrasl_0(xrasl[0]),
	.xrasl_1(xrasl[1]),
	.xdtackl(xdtackl),
	.xintl(xintl),
	.hs_o(hs_o),
	.hhs_o(hhs_o),
	.vs_o(vs_o),
	.refreq(refreq),
	.obbreq(obbreq),
	.bbreq_0(bbreq[0]),
	.bbreq_1(bbreq[1]),
	.gbreq_0(gbreq[0]),
	.gbreq_1(gbreq[1]),
	.dram(fdram),	// /!\
	.blank(blank),
	.tlw(tlw),
	.ram_rdy(ram_rdy),
	.aen(aen),
	.den_0(den[0]),
	.den_1(den[1]),
	.den_2(den[2]),
	.sys_clk(sys_clk),
	.startcas(startcas),
	.hsl(hsl),
	.vsl(vsl)
);

endmodule
