module j_jbus
(
	input ain_0,
	input ain_1,
	input ain_2,
	input ain_3,
	input ain_4,
	input ain_5,
	input ain_6,
	input ain_7,
	input ain_8,
	input ain_9,
	input ain_10,
	input ain_11,
	input ain_12,
	input ain_13,
	input ain_14,
	input ain_15,
	input ain_16,
	input ain_17,
	input ain_18,
	input ain_19,
	input ain_20,
	input ain_21,
	input ain_22,
	input ain_23,
	input din_0,
	input din_1,
	input din_2,
	input din_3,
	input din_4,
	input din_5,
	input din_6,
	input din_7,
	input din_8,
	input din_9,
	input din_10,
	input din_11,
	input din_12,
	input din_13,
	input din_14,
	input din_15,
	input din_16,
	input din_17,
	input din_18,
	input din_19,
	input din_20,
	input din_21,
	input din_22,
	input din_23,
	input din_24,
	input din_25,
	input din_26,
	input din_27,
	input din_28,
	input din_29,
	input din_30,
	input din_31,
	input dr_0,
	input dr_1,
	input dr_2,
	input dr_3,
	input dr_4,
	input dr_5,
	input dr_6,
	input dr_7,
	input dr_8,
	input dr_9,
	input dr_10,
	input dr_11,
	input dr_12,
	input dr_13,
	input dr_14,
	input dr_15,
	input dinlatch_0,
	input dinlatch_1,
	input dmuxd_0,
	input dmuxd_1,
	input dmuxu_0,
	input dmuxu_1,
	input dren,
	input xdsrc,
	input ack,
	input wd_0,
	input wd_1,
	input wd_2,
	input wd_3,
	input wd_4,
	input wd_5,
	input wd_6,
	input wd_7,
	input wd_8,
	input wd_9,
	input wd_10,
	input wd_11,
	input wd_12,
	input wd_13,
	input wd_14,
	input wd_15,
	input wd_16,
	input wd_17,
	input wd_18,
	input wd_19,
	input wd_20,
	input wd_21,
	input wd_22,
	input wd_23,
	input wd_24,
	input wd_25,
	input wd_26,
	input wd_27,
	input wd_28,
	input wd_29,
	input wd_30,
	input wd_31,
	input clk,
	input cfg_0,
	input cfg_1,
	input cfgw,
	input a_0,
	input a_1,
	input a_2,
	input a_3,
	input a_4,
	input a_5,
	input a_6,
	input a_7,
	input a_8,
	input a_9,
	input a_10,
	input a_11,
	input a_12,
	input a_13,
	input a_14,
	input a_15,
	input a_16,
	input a_17,
	input a_18,
	input a_19,
	input a_20,
	input a_21,
	input a_22,
	input a_23,
	input ainen,
	input seta1,
	input masterdata,
	output dout_0,
	output dout_1,
	output dout_2,
	output dout_3,
	output dout_4,
	output dout_5,
	output dout_6,
	output dout_7,
	output dout_8,
	output dout_9,
	output dout_10,
	output dout_11,
	output dout_12,
	output dout_13,
	output dout_14,
	output dout_15,
	output dout_16,
	output dout_17,
	output dout_18,
	output dout_19,
	output dout_20,
	output dout_21,
	output dout_22,
	output dout_23,
	output dout_24,
	output dout_25,
	output dout_26,
	output dout_27,
	output dout_28,
	output dout_29,
	output dout_30,
	output dout_31,
	output aout_0,
	output aout_1,
	output aout_2,
	output aout_3,
	output aout_4,
	output aout_5,
	output aout_6,
	output aout_7,
	output aout_8,
	output aout_9,
	output aout_10,
	output aout_11,
	output aout_12,
	output aout_13,
	output aout_14,
	output aout_15,
	output aout_16,
	output aout_17,
	output aout_18,
	output aout_19,
	output aout_20,
	output aout_21,
	output aout_22,
	output aout_23,
	output dsp16,
	output bigend,
	input sys_clk // Generated
);
wire [23:0] ain = {ain_23,ain_22,ain_21,ain_20,
ain_19,ain_18,ain_17,ain_16,ain_15,ain_14,ain_13,ain_12,ain_11,ain_10,
ain_9,ain_8,ain_7,ain_6,ain_5,ain_4,ain_3,ain_2,ain_1,ain_0};
wire [31:0] din = {din_31,din_30,
din_29,din_28,din_27,din_26,din_25,din_24,din_23,din_22,din_21,din_20,
din_19,din_18,din_17,din_16,din_15,din_14,din_13,din_12,din_11,din_10,
din_9,din_8,din_7,din_6,din_5,din_4,din_3,din_2,din_1,din_0};
wire [15:0] dr = {dr_15,dr_14,dr_13,dr_12,dr_11,dr_10,
dr_9,dr_8,dr_7,dr_6,dr_5,dr_4,dr_3,dr_2,dr_1,dr_0};
wire [1:0] dinlatch = {dinlatch_1,dinlatch_0};
wire [1:0] dmuxd = {dmuxd_1,dmuxd_0};
wire [1:0] dmuxu = {dmuxu_1,dmuxu_0};
wire [31:0] wd = {wd_31,wd_30,
wd_29,wd_28,wd_27,wd_26,wd_25,wd_24,wd_23,wd_22,wd_21,wd_20,
wd_19,wd_18,wd_17,wd_16,wd_15,wd_14,wd_13,wd_12,wd_11,wd_10,
wd_9,wd_8,wd_7,wd_6,wd_5,wd_4,wd_3,wd_2,wd_1,wd_0};
wire [1:0] cfg = {cfg_1,cfg_0};
wire [23:0] a = {a_23,a_22,a_21,a_20,
a_19,a_18,a_17,a_16,a_15,a_14,a_13,a_12,a_11,a_10,
a_9,a_8,a_7,a_6,a_5,a_4,a_3,a_2,a_1,a_0};
wire [31:0] dout;
assign {dout_31,dout_30,
dout_29,dout_28,dout_27,dout_26,dout_25,dout_24,dout_23,dout_22,dout_21,dout_20,
dout_19,dout_18,dout_17,dout_16,dout_15,dout_14,dout_13,dout_12,dout_11,dout_10,
dout_9,dout_8,dout_7,dout_6,dout_5,dout_4,dout_3,dout_2,dout_1,dout_0} = dout[31:0];
wire [23:0] aout;
assign {aout_23,aout_22,aout_21,aout_20,
aout_19,aout_18,aout_17,aout_16,aout_15,aout_14,aout_13,aout_12,aout_11,aout_10,
aout_9,aout_8,aout_7,aout_6,aout_5,aout_4,aout_3,aout_2,aout_1,aout_0} = aout[23:0];
_j_jbus jbus_inst
(
	.ain /* IN */ (ain[23:0]),
	.din /* IN */ (din[31:0]),
	.dr /* IN */ (dr[15:0]),
	.dinlatch /* IN */ (dinlatch[1:0]),
	.dmuxd /* IN */ (dmuxd[1:0]),
	.dmuxu /* IN */ (dmuxu[1:0]),
	.dren /* IN */ (dren),
	.xdsrc /* IN */ (xdsrc),
	.ack /* IN */ (ack),
	.wd /* IN */ (wd[31:0]),
	.clk /* IN */ (clk),
	.cfg /* IN */ (cfg[1:0]),
	.cfgw /* IN */ (cfgw),
	.a /* IN */ (a[23:0]),
	.ainen /* IN */ (ainen),
	.seta1 /* IN */ (seta1),
	.masterdata /* IN */ (masterdata),
	.dout /* OUT */ (dout[31:0]),
	.aout /* OUT */ (aout[23:0]),
	.dsp16 /* OUT */ (dsp16),
	.bigend /* OUT */ (bigend),
	.sys_clk(sys_clk) // Generated
);
endmodule
