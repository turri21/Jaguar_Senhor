module data
(
	output wdata_0_out,
	output wdata_0_oe,
	input wdata_0_in,
	output wdata_1_out,
	output wdata_1_oe,
	input wdata_1_in,
	output wdata_2_out,
	output wdata_2_oe,
	input wdata_2_in,
	output wdata_3_out,
	output wdata_3_oe,
	input wdata_3_in,
	output wdata_4_out,
	output wdata_4_oe,
	input wdata_4_in,
	output wdata_5_out,
	output wdata_5_oe,
	input wdata_5_in,
	output wdata_6_out,
	output wdata_6_oe,
	input wdata_6_in,
	output wdata_7_out,
	output wdata_7_oe,
	input wdata_7_in,
	output wdata_8_out,
	output wdata_8_oe,
	input wdata_8_in,
	output wdata_9_out,
	output wdata_9_oe,
	input wdata_9_in,
	output wdata_10_out,
	output wdata_10_oe,
	input wdata_10_in,
	output wdata_11_out,
	output wdata_11_oe,
	input wdata_11_in,
	output wdata_12_out,
	output wdata_12_oe,
	input wdata_12_in,
	output wdata_13_out,
	output wdata_13_oe,
	input wdata_13_in,
	output wdata_14_out,
	output wdata_14_oe,
	input wdata_14_in,
	output wdata_15_out,
	output wdata_15_oe,
	input wdata_15_in,
	output wdata_16_out,
	output wdata_16_oe,
	input wdata_16_in,
	output wdata_17_out,
	output wdata_17_oe,
	input wdata_17_in,
	output wdata_18_out,
	output wdata_18_oe,
	input wdata_18_in,
	output wdata_19_out,
	output wdata_19_oe,
	input wdata_19_in,
	output wdata_20_out,
	output wdata_20_oe,
	input wdata_20_in,
	output wdata_21_out,
	output wdata_21_oe,
	input wdata_21_in,
	output wdata_22_out,
	output wdata_22_oe,
	input wdata_22_in,
	output wdata_23_out,
	output wdata_23_oe,
	input wdata_23_in,
	output wdata_24_out,
	output wdata_24_oe,
	input wdata_24_in,
	output wdata_25_out,
	output wdata_25_oe,
	input wdata_25_in,
	output wdata_26_out,
	output wdata_26_oe,
	input wdata_26_in,
	output wdata_27_out,
	output wdata_27_oe,
	input wdata_27_in,
	output wdata_28_out,
	output wdata_28_oe,
	input wdata_28_in,
	output wdata_29_out,
	output wdata_29_oe,
	input wdata_29_in,
	output wdata_30_out,
	output wdata_30_oe,
	input wdata_30_in,
	output wdata_31_out,
	output wdata_31_oe,
	input wdata_31_in,
	output wdata_32_out,
	output wdata_32_oe,
	input wdata_32_in,
	output wdata_33_out,
	output wdata_33_oe,
	input wdata_33_in,
	output wdata_34_out,
	output wdata_34_oe,
	input wdata_34_in,
	output wdata_35_out,
	output wdata_35_oe,
	input wdata_35_in,
	output wdata_36_out,
	output wdata_36_oe,
	input wdata_36_in,
	output wdata_37_out,
	output wdata_37_oe,
	input wdata_37_in,
	output wdata_38_out,
	output wdata_38_oe,
	input wdata_38_in,
	output wdata_39_out,
	output wdata_39_oe,
	input wdata_39_in,
	output wdata_40_out,
	output wdata_40_oe,
	input wdata_40_in,
	output wdata_41_out,
	output wdata_41_oe,
	input wdata_41_in,
	output wdata_42_out,
	output wdata_42_oe,
	input wdata_42_in,
	output wdata_43_out,
	output wdata_43_oe,
	input wdata_43_in,
	output wdata_44_out,
	output wdata_44_oe,
	input wdata_44_in,
	output wdata_45_out,
	output wdata_45_oe,
	input wdata_45_in,
	output wdata_46_out,
	output wdata_46_oe,
	input wdata_46_in,
	output wdata_47_out,
	output wdata_47_oe,
	input wdata_47_in,
	output wdata_48_out,
	output wdata_48_oe,
	input wdata_48_in,
	output wdata_49_out,
	output wdata_49_oe,
	input wdata_49_in,
	output wdata_50_out,
	output wdata_50_oe,
	input wdata_50_in,
	output wdata_51_out,
	output wdata_51_oe,
	input wdata_51_in,
	output wdata_52_out,
	output wdata_52_oe,
	input wdata_52_in,
	output wdata_53_out,
	output wdata_53_oe,
	input wdata_53_in,
	output wdata_54_out,
	output wdata_54_oe,
	input wdata_54_in,
	output wdata_55_out,
	output wdata_55_oe,
	input wdata_55_in,
	output wdata_56_out,
	output wdata_56_oe,
	input wdata_56_in,
	output wdata_57_out,
	output wdata_57_oe,
	input wdata_57_in,
	output wdata_58_out,
	output wdata_58_oe,
	input wdata_58_in,
	output wdata_59_out,
	output wdata_59_oe,
	input wdata_59_in,
	output wdata_60_out,
	output wdata_60_oe,
	input wdata_60_in,
	output wdata_61_out,
	output wdata_61_oe,
	input wdata_61_in,
	output wdata_62_out,
	output wdata_62_oe,
	input wdata_62_in,
	output wdata_63_out,
	output wdata_63_oe,
	input wdata_63_in,
	output dcomp_0,
	output dcomp_1,
	output dcomp_2,
	output dcomp_3,
	output dcomp_4,
	output dcomp_5,
	output dcomp_6,
	output dcomp_7,
	output srcd_0,
	output srcd_1,
	output srcd_2,
	output srcd_3,
	output srcd_4,
	output srcd_5,
	output srcd_6,
	output srcd_7,
	output zcomp_0,
	output zcomp_1,
	output zcomp_2,
	output zcomp_3,
	input big_pix,
	input blit_back,
	input blit_breq_0,
	input blit_breq_1,
	input clk,
	input clk2,
	input cmpdst,
	input daddasel_0,
	input daddasel_1,
	input daddasel_2,
	input daddbsel_0,
	input daddbsel_1,
	input daddbsel_2,
	input daddmode_0,
	input daddmode_1,
	input daddmode_2,
	input daddq_sel,
	input data_0,
	input data_1,
	input data_2,
	input data_3,
	input data_4,
	input data_5,
	input data_6,
	input data_7,
	input data_8,
	input data_9,
	input data_10,
	input data_11,
	input data_12,
	input data_13,
	input data_14,
	input data_15,
	input data_16,
	input data_17,
	input data_18,
	input data_19,
	input data_20,
	input data_21,
	input data_22,
	input data_23,
	input data_24,
	input data_25,
	input data_26,
	input data_27,
	input data_28,
	input data_29,
	input data_30,
	input data_31,
	input data_32,
	input data_33,
	input data_34,
	input data_35,
	input data_36,
	input data_37,
	input data_38,
	input data_39,
	input data_40,
	input data_41,
	input data_42,
	input data_43,
	input data_44,
	input data_45,
	input data_46,
	input data_47,
	input data_48,
	input data_49,
	input data_50,
	input data_51,
	input data_52,
	input data_53,
	input data_54,
	input data_55,
	input data_56,
	input data_57,
	input data_58,
	input data_59,
	input data_60,
	input data_61,
	input data_62,
	input data_63,
	input data_ena,
	input data_sel_0,
	input data_sel_1,
	input dbinh_n_0,
	input dbinh_n_1,
	input dbinh_n_2,
	input dbinh_n_3,
	input dbinh_n_4,
	input dbinh_n_5,
	input dbinh_n_6,
	input dbinh_n_7,
	input dend_0,
	input dend_1,
	input dend_2,
	input dend_3,
	input dend_4,
	input dend_5,
	input dpipe_0,
	input dpipe_1,
	input dstart_0,
	input dstart_1,
	input dstart_2,
	input dstart_3,
	input dstart_4,
	input dstart_5,
	input dstdld_0,
	input dstdld_1,
	input dstzld_0,
	input dstzld_1,
	input [0:31] gpu_din,
	input iincld,
	input intld_0,
	input intld_1,
	input intld_2,
	input intld_3,
	input lfu_func_0,
	input lfu_func_1,
	input lfu_func_2,
	input lfu_func_3,
	input load_strobe,
	input patdld_0,
	input patdld_1,
	input phrase_mode,
	input reset_n,
	input srcd1ld_0,
	input srcd1ld_1,
	input srcdread,
	input srczread,
	input srcshift_0,
	input srcshift_1,
	input srcshift_2,
	input srcshift_3,
	input srcshift_4,
	input srcshift_5,
	input srcz1ld_0,
	input srcz1ld_1,
	input srcz2add,
	input srcz2ld_0,
	input srcz2ld_1,
	input zedld_0,
	input zedld_1,
	input zedld_2,
	input zedld_3,
	input zincld,
	input zmode_0,
	input zmode_1,
	input zmode_2,
	input zpipe_0,
	input zpipe_1,
	input sys_clk // Generated
);
wire [63:0] wdata_out;
assign {wdata_63_out,wdata_62_out,wdata_61_out,wdata_60_out,
wdata_59_out,wdata_58_out,wdata_57_out,wdata_56_out,wdata_55_out,wdata_54_out,wdata_53_out,wdata_52_out,wdata_51_out,wdata_50_out,
wdata_49_out,wdata_48_out,wdata_47_out,wdata_46_out,wdata_45_out,wdata_44_out,wdata_43_out,wdata_42_out,wdata_41_out,wdata_40_out,
wdata_39_out,wdata_38_out,wdata_37_out,wdata_36_out,wdata_35_out,wdata_34_out,wdata_33_out,wdata_32_out,wdata_31_out,wdata_30_out,
wdata_29_out,wdata_28_out,wdata_27_out,wdata_26_out,wdata_25_out,wdata_24_out,wdata_23_out,wdata_22_out,wdata_21_out,wdata_20_out,
wdata_19_out,wdata_18_out,wdata_17_out,wdata_16_out,wdata_15_out,wdata_14_out,wdata_13_out,wdata_12_out,wdata_11_out,wdata_10_out,
wdata_9_out,wdata_8_out,wdata_7_out,wdata_6_out,wdata_5_out,wdata_4_out,wdata_3_out,wdata_2_out,wdata_1_out,wdata_0_out} = wdata_out[63:0];
assign {wdata_63_oe,wdata_62_oe,wdata_61_oe,wdata_60_oe,
wdata_59_oe,wdata_58_oe,wdata_57_oe,wdata_56_oe,wdata_55_oe,wdata_54_oe,wdata_53_oe,wdata_52_oe,wdata_51_oe,wdata_50_oe,
wdata_49_oe,wdata_48_oe,wdata_47_oe,wdata_46_oe,wdata_45_oe,wdata_44_oe,wdata_43_oe,wdata_42_oe,wdata_41_oe,wdata_40_oe,
wdata_39_oe,wdata_38_oe,wdata_37_oe,wdata_36_oe,wdata_35_oe,wdata_34_oe,wdata_33_oe,wdata_32_oe,wdata_31_oe,wdata_30_oe,
wdata_29_oe,wdata_28_oe,wdata_27_oe,wdata_26_oe,wdata_25_oe,wdata_24_oe,wdata_23_oe,wdata_22_oe,wdata_21_oe,wdata_20_oe,
wdata_19_oe,wdata_18_oe,wdata_17_oe,wdata_16_oe,wdata_15_oe,wdata_14_oe,wdata_13_oe,wdata_12_oe,wdata_11_oe,wdata_10_oe,
wdata_9_oe,wdata_8_oe,wdata_7_oe,wdata_6_oe,wdata_5_oe,wdata_4_oe,wdata_3_oe,wdata_2_oe,wdata_1_oe} = {63{wdata_0_oe}};
wire [7:0] dcomp;
assign {dcomp_7,dcomp_6,dcomp_5,dcomp_4,dcomp_3,dcomp_2,dcomp_1,dcomp_0} = dcomp[7:0];
wire [7:0] srcd;
assign {srcd_7,srcd_6,srcd_5,srcd_4,srcd_3,srcd_2,srcd_1,srcd_0} = srcd[7:0];
wire [3:0] zcomp;
assign {zcomp_3,zcomp_2,zcomp_1,zcomp_0} = zcomp[3:0];
wire [1:0] blit_breq = {blit_breq_1,blit_breq_0};
wire [2:0] daddasel = {daddasel_2,daddasel_1,daddasel_0};
wire [2:0] daddbsel = {daddbsel_2,daddbsel_1,daddbsel_0};
wire [2:0] daddmode = {daddmode_2,daddmode_1,daddmode_0};
wire [63:0] data = {data_63,data_62,data_61,data_60,
data_59,data_58,data_57,data_56,data_55,data_54,data_53,data_52,data_51,data_50,
data_49,data_48,data_47,data_46,data_45,data_44,data_43,data_42,data_41,data_40,
data_39,data_38,data_37,data_36,data_35,data_34,data_33,data_32,data_31,data_30,
data_29,data_28,data_27,data_26,data_25,data_24,data_23,data_22,data_21,data_20,
data_19,data_18,data_17,data_16,data_15,data_14,data_13,data_12,data_11,data_10,
data_9,data_8,data_7,data_6,data_5,data_4,data_3,data_2,data_1,data_0};
wire [1:0] data_sel = {data_sel_1,data_sel_0};
wire [7:0] dbinh_n = {dbinh_n_7,dbinh_n_6,dbinh_n_5,dbinh_n_4,dbinh_n_3,dbinh_n_2,dbinh_n_1,dbinh_n_0};
wire [5:0] dend = {dend_5,dend_4,dend_3,dend_2,dend_1,dend_0};
wire [1:0] dpipe = {dpipe_1,dpipe_0};
wire [5:0] dstart = {dstart_5,dstart_4,dstart_3,dstart_2,dstart_1,dstart_0};
wire [1:0] dstdld = {dstdld_1,dstdld_0};
wire [1:0] dstzld = {dstzld_1,dstzld_0};
wire [31:0] gpu_din_ = {gpu_din[31],gpu_din[30],
gpu_din[29],gpu_din[28],gpu_din[27],gpu_din[26],gpu_din[25],gpu_din[24],gpu_din[23],gpu_din[22],gpu_din[21],gpu_din[20],
gpu_din[19],gpu_din[18],gpu_din[17],gpu_din[16],gpu_din[15],gpu_din[14],gpu_din[13],gpu_din[12],gpu_din[11],gpu_din[10],
gpu_din[9],gpu_din[8],gpu_din[7],gpu_din[6],gpu_din[5],gpu_din[4],gpu_din[3],gpu_din[2],gpu_din[1],gpu_din[0]};
wire [3:0] intld = {intld_3,intld_2,intld_1,intld_0};
wire [3:0] lfu_func = {lfu_func_3,lfu_func_2,lfu_func_1,lfu_func_0};
wire [1:0] patdld = {patdld_1,patdld_0};
wire [1:0] srcd1ld = {srcd1ld_1,srcd1ld_0};
wire [5:0] srcshift = {srcshift_5,srcshift_4,srcshift_3,srcshift_2,srcshift_1,srcshift_0};
wire [1:0] srcz1ld = {srcz1ld_1,srcz1ld_0};
wire [1:0] srcz2ld = {srcz2ld_1,srcz2ld_0};
wire [3:0] zedld = {zedld_3,zedld_2,zedld_1,zedld_0};
wire [2:0] zmode = {zmode_2,zmode_1,zmode_0};
wire [1:0] zpipe = {zpipe_1,zpipe_0};

_data data_inst
(
	.wdata_out /* BUS */ (wdata_out[63:0]),
	.wdata_oe /* BUS */ (wdata_0_oe),
	.dcomp /* OUT */ (dcomp[7:0]),
	.srcd /* OUT */ (srcd[7:0]),
	.zcomp /* OUT */ (zcomp[3:0]),
	.big_pix /* IN */ (big_pix),
	.blit_back /* IN */ (blit_back),
	.blit_breq /* IN */ (blit_breq[1:0]),
	.clk /* IN */ (clk),
	.clk2 /* IN */ (clk2),
	.cmpdst /* IN */ (cmpdst),
	.daddasel /* IN */ (daddasel[2:0]),
	.daddbsel /* IN */ (daddbsel[2:0]),
	.daddmode /* IN */ (daddmode[2:0]),
	.daddq_sel /* IN */ (daddq_sel),
	.data /* IN */ (data[63:0]),
	.data_ena /* IN */ (data_ena),
	.data_sel /* IN */ (data_sel[1:0]),
	.dbinh_n /* IN */ (dbinh_n[7:0]),
	.dend /* IN */ (dend[5:0]),
	.dpipe /* IN */ (dpipe[1:0]),
	.dstart /* IN */ (dstart[5:0]),
	.dstdld /* IN */ (dstdld[1:0]),
	.dstzld /* IN */ (dstzld[1:0]),
	.gpu_din /* IN */ (gpu_din_[31:0]),
	.iincld /* IN */ (iincld),
	.intld /* IN */ (intld[3:0]),
	.lfu_func /* IN */ (lfu_func[3:0]),
	.load_strobe /* IN */ (load_strobe),
	.patdld /* IN */ (patdld[1:0]),
	.phrase_mode /* IN */ (phrase_mode),
	.reset_n /* IN */ (reset_n),
	.srcd1ld /* IN */ (srcd1ld[1:0]),
	.srcdread /* IN */ (srcdread),
	.srczread /* IN */ (srczread),
	.srcshift /* IN */ (srcshift[5:0]),
	.srcz1ld /* IN */ (srcz1ld[1:0]),
	.srcz2add /* IN */ (srcz2add),
	.srcz2ld /* IN */ (srcz2ld[1:0]),
	.zedld /* IN */ (zedld[3:0]),
	.zincld /* IN */ (zincld),
	.zmode /* IN */ (zmode[2:0]),
	.zpipe /* IN */ (zpipe[1:0]),
	.sys_clk(sys_clk) // Generated
);
endmodule
