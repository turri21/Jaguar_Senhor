module state
(
	output [0:23] blit_addr_out,
	output blit_addr_oe,
	input [0:23] blit_addr_in,
	output justify_out,
	output justify_oe,
	input justify_in,
	output mreq_out,
	output mreq_oe,
	input mreq_in,
	output width_0_out,
	output width_0_oe,
	input width_0_in,
	output width_1_out,
	output width_1_oe,
	input width_1_in,
	output width_2_out,
	output width_2_oe,
	input width_2_in,
	output width_3_out,
	output width_3_oe,
	input width_3_in,
	output read_out,
	output read_oe,
	input read_in,
	output gpu_dout_0_out,
	output gpu_dout_0_oe,
	input gpu_dout_0_in,
	output gpu_dout_1_out,
	output gpu_dout_1_oe,
	input gpu_dout_1_in,
	output gpu_dout_2_out,
	output gpu_dout_2_oe,
	input gpu_dout_2_in,
	output gpu_dout_3_out,
	output gpu_dout_3_oe,
	input gpu_dout_3_in,
	output gpu_dout_4_out,
	output gpu_dout_4_oe,
	input gpu_dout_4_in,
	output gpu_dout_5_out,
	output gpu_dout_5_oe,
	input gpu_dout_5_in,
	output gpu_dout_6_out,
	output gpu_dout_6_oe,
	input gpu_dout_6_in,
	output gpu_dout_7_out,
	output gpu_dout_7_oe,
	input gpu_dout_7_in,
	output gpu_dout_8_out,
	output gpu_dout_8_oe,
	input gpu_dout_8_in,
	output gpu_dout_9_out,
	output gpu_dout_9_oe,
	input gpu_dout_9_in,
	output gpu_dout_10_out,
	output gpu_dout_10_oe,
	input gpu_dout_10_in,
	output gpu_dout_11_out,
	output gpu_dout_11_oe,
	input gpu_dout_11_in,
	output gpu_dout_12_out,
	output gpu_dout_12_oe,
	input gpu_dout_12_in,
	output gpu_dout_13_out,
	output gpu_dout_13_oe,
	input gpu_dout_13_in,
	output gpu_dout_14_out,
	output gpu_dout_14_oe,
	input gpu_dout_14_in,
	output gpu_dout_15_out,
	output gpu_dout_15_oe,
	input gpu_dout_15_in,
	output gpu_dout_16_out,
	output gpu_dout_16_oe,
	input gpu_dout_16_in,
	output gpu_dout_17_out,
	output gpu_dout_17_oe,
	input gpu_dout_17_in,
	output gpu_dout_18_out,
	output gpu_dout_18_oe,
	input gpu_dout_18_in,
	output gpu_dout_19_out,
	output gpu_dout_19_oe,
	input gpu_dout_19_in,
	output gpu_dout_20_out,
	output gpu_dout_20_oe,
	input gpu_dout_20_in,
	output gpu_dout_21_out,
	output gpu_dout_21_oe,
	input gpu_dout_21_in,
	output gpu_dout_22_out,
	output gpu_dout_22_oe,
	input gpu_dout_22_in,
	output gpu_dout_23_out,
	output gpu_dout_23_oe,
	input gpu_dout_23_in,
	output gpu_dout_24_out,
	output gpu_dout_24_oe,
	input gpu_dout_24_in,
	output gpu_dout_25_out,
	output gpu_dout_25_oe,
	input gpu_dout_25_in,
	output gpu_dout_26_out,
	output gpu_dout_26_oe,
	input gpu_dout_26_in,
	output gpu_dout_27_out,
	output gpu_dout_27_oe,
	input gpu_dout_27_in,
	output gpu_dout_28_out,
	output gpu_dout_28_oe,
	input gpu_dout_28_in,
	output gpu_dout_29_out,
	output gpu_dout_29_oe,
	input gpu_dout_29_in,
	output gpu_dout_30_out,
	output gpu_dout_30_oe,
	input gpu_dout_30_in,
	output gpu_dout_31_out,
	output gpu_dout_31_oe,
	input gpu_dout_31_in,
	output a1fracldi,
	output a1ptrldi,
	output a2ptrldi,
	output addasel_0,
	output addasel_1,
	output addasel_2,
	output addbsel_0,
	output addbsel_1,
	output addqsel,
	output adda_xconst_0,
	output adda_xconst_1,
	output adda_xconst_2,
	output adda_yconst,
	output addareg,
	output apipe,
	output blit_breq_0,
	output blit_breq_1,
	output blit_int,
	output cmpdst,
	output daddasel_0,
	output daddasel_1,
	output daddasel_2,
	output daddbsel_0,
	output daddbsel_1,
	output daddbsel_2,
	output daddmode_0,
	output daddmode_1,
	output daddmode_2,
	output data_ena,
	output data_sel_0,
	output data_sel_1,
	output dbinh_n_0,
	output dbinh_n_1,
	output dbinh_n_2,
	output dbinh_n_3,
	output dbinh_n_4,
	output dbinh_n_5,
	output dbinh_n_6,
	output dbinh_n_7,
	output dend_0,
	output dend_1,
	output dend_2,
	output dend_3,
	output dend_4,
	output dend_5,
	output dpipe_0,
	output dpipe_1,
	output dstart_0,
	output dstart_1,
	output dstart_2,
	output dstart_3,
	output dstart_4,
	output dstart_5,
	output dstdread,
	output dstzread,
	output gena2,
	output lfu_func_0,
	output lfu_func_1,
	output lfu_func_2,
	output lfu_func_3,
	output daddq_sel,
	output modx_0,
	output modx_1,
	output modx_2,
	output patdadd,
	output patfadd,
	output phrase_mode,
	output reset_n,
	output srcdread,
	output srcshift_0,
	output srcshift_1,
	output srcshift_2,
	output srcshift_3,
	output srcshift_4,
	output srcshift_5,
	output srcz1add,
	output srcz2add,
	output srczread,
	output suba_x,
	output suba_y,
	output zaddr,
	output zmode_0,
	output zmode_1,
	output zmode_2,
	output zpipe_0,
	output zpipe_1,
	input a1_outside,
	input a1_pixsize_0,
	input a1_pixsize_1,
	input a1_pixsize_2,
	input [0:14] a1_win_x,
	input [0:15] a1_x,
	input a1addx_0,
	input a1addx_1,
	input a1addy,
	input a1xsign,
	input a1ysign,
	input a2_pixsize_0,
	input a2_pixsize_1,
	input a2_pixsize_2,
	input [0:15] a2_x,
	input a2addx_0,
	input a2addx_1,
	input a2addy,
	input a2xsign,
	input a2ysign,
	input ack,
	input [0:23] address,
	input big_pix,
	input blit_back,
	input clk,
	input cmdld,
	input countld,
	input dcomp_0,
	input dcomp_1,
	input dcomp_2,
	input dcomp_3,
	input dcomp_4,
	input dcomp_5,
	input dcomp_6,
	input dcomp_7,
	input [0:31] gpu_din,
	input pixa_0,
	input pixa_1,
	input pixa_2,
	input srcd_0,
	input srcd_1,
	input srcd_2,
	input srcd_3,
	input srcd_4,
	input srcd_5,
	input srcd_6,
	input srcd_7,
	input statrd,
	input stopld,
	input xreset_n,
	input zcomp_0,
	input zcomp_1,
	input zcomp_2,
	input zcomp_3,
	input sys_clk // Generated
);

wire [23:0] blit_addr_out_;
assign {blit_addr_out[23],blit_addr_out[22],blit_addr_out[21],blit_addr_out[20],
blit_addr_out[19],blit_addr_out[18],blit_addr_out[17],blit_addr_out[16],blit_addr_out[15],blit_addr_out[14],blit_addr_out[13],blit_addr_out[12],blit_addr_out[11],blit_addr_out[10],
blit_addr_out[9],blit_addr_out[8],blit_addr_out[7],blit_addr_out[6],blit_addr_out[5],blit_addr_out[4],blit_addr_out[3],blit_addr_out[2],blit_addr_out[1],blit_addr_out[0]} = blit_addr_out_[23:0];
wire [3:0] width_out;
assign {width_3_out,width_2_out,width_1_out,width_0_out} = width_out[3:0];
assign {width_3_oe,width_2_oe,width_1_oe} = {3{width_0_oe}};
wire [31:0] gpu_dout_out;
assign {gpu_dout_31_out,gpu_dout_30_out,
gpu_dout_29_out,gpu_dout_28_out,gpu_dout_27_out,gpu_dout_26_out,gpu_dout_25_out,gpu_dout_24_out,gpu_dout_23_out,gpu_dout_22_out,gpu_dout_21_out,gpu_dout_20_out,
gpu_dout_19_out,gpu_dout_18_out,gpu_dout_17_out,gpu_dout_16_out,gpu_dout_15_out,gpu_dout_14_out,gpu_dout_13_out,gpu_dout_12_out,gpu_dout_11_out,gpu_dout_10_out,
gpu_dout_9_out,gpu_dout_8_out,gpu_dout_7_out,gpu_dout_6_out,gpu_dout_5_out,gpu_dout_4_out,gpu_dout_3_out,gpu_dout_2_out,gpu_dout_1_out,gpu_dout_0_out,} = gpu_dout_out[31:0];
assign {gpu_dout_31_oe,gpu_dout_30_oe,
gpu_dout_29_oe,gpu_dout_28_oe,gpu_dout_27_oe,gpu_dout_26_oe,gpu_dout_25_oe,gpu_dout_24_oe,gpu_dout_23_oe,gpu_dout_22_oe,gpu_dout_21_oe,gpu_dout_20_oe,
gpu_dout_19_oe,gpu_dout_18_oe,gpu_dout_17_oe,gpu_dout_16_oe,gpu_dout_15_oe,gpu_dout_14_oe,gpu_dout_13_oe,gpu_dout_12_oe,gpu_dout_11_oe,gpu_dout_10_oe,
gpu_dout_9_oe,gpu_dout_8_oe,gpu_dout_7_oe,gpu_dout_6_oe,gpu_dout_5_oe,gpu_dout_4_oe,gpu_dout_3_oe,gpu_dout_2_oe,gpu_dout_1_oe,gpu_dout_0_oe,} = {31{gpu_dout_0_oe}};
wire [2:0] addasel;
assign {addasel_2,addasel_1,addasel_0} = addasel[2:0];
wire [1:0] addbsel;
assign {addbsel_1,addbsel_0} = addbsel[1:0];
wire [2:0] adda_xconst;
assign {adda_xconst_2,adda_xconst_1,adda_xconst_0} = adda_xconst[2:0];
wire [1:0] blit_breq;
assign {blit_breq_1,blit_breq_0} = blit_breq[1:0];
wire [2:0] daddasel;
assign {daddasel_2,daddasel_1,daddasel_0} = daddasel[2:0];
wire [2:0] daddbsel;
assign {daddbsel_2,daddbsel_1,daddbsel_0} = daddbsel[2:0];
wire [2:0] daddmode;
assign {daddmode_2,daddmode_1,daddmode_0} = daddmode[2:0];
wire [1:0] data_sel;
assign {data_sel_1,data_sel_0} = data_sel[1:0];
wire [7:0] dbinh_n;
assign {dbinh_n_7,dbinh_n_6,dbinh_n_5,dbinh_n_4,dbinh_n_3,dbinh_n_2,dbinh_n_1,dbinh_n_0} = dbinh_n[7:0];
wire [5:0] dend;
assign {dend_5,dend_4,dend_3,dend_2,dend_1,dend_0} = dend[5:0];
wire [1:0] dpipe;
assign {dpipe_1,dpipe_0} = dpipe[1:0];
wire [5:0] dstart;
assign {dstart_5,dstart_4,dstart_3,dstart_2,dstart_1,dstart_0} = dstart[5:0];
wire [3:0] lfu_func;
assign {lfu_func_3,lfu_func_2,lfu_func_1,lfu_func_0} = lfu_func[3:0];
wire [2:0] modx;
assign {modx_2,modx_1,modx_0} = modx[2:0];
wire [5:0] srcshift;
assign {srcshift_5,srcshift_4,srcshift_3,srcshift_2,srcshift_1,srcshift_0} = srcshift[5:0];
wire [2:0] zmode;
assign {zmode_2,zmode_1,zmode_0} = zmode[2:0];
wire [1:0] zpipe;
assign {zpipe_1,zpipe_0} = zpipe[1:0];
wire [2:0] a1_pixsize = {a1_pixsize_2,a1_pixsize_1,a1_pixsize_0};
wire [14:0] a1_win_x_ = {a1_win_x[14],a1_win_x[13],a1_win_x[12],a1_win_x[11],a1_win_x[10],
a1_win_x[9],a1_win_x[8],a1_win_x[7],a1_win_x[6],a1_win_x[5],a1_win_x[4],a1_win_x[3],a1_win_x[2],a1_win_x[1],a1_win_x[0]};
wire [15:0] a1_x_ = {a1_x[15],a1_x[14],a1_x[13],a1_x[12],a1_x[11],a1_x[10],
a1_x[9],a1_x[8],a1_x[7],a1_x[6],a1_x[5],a1_x[4],a1_x[3],a1_x[2],a1_x[1],a1_x[0]};
wire [1:0] a1addx = {a1addx_1,a1addx_0};
wire [2:0] a2_pixsize = {a2_pixsize_2,a2_pixsize_1,a2_pixsize_0};
wire [15:0] a2_x_ = {a2_x[15],a2_x[14],a2_x[13],a2_x[12],a2_x[11],a2_x[10],
a2_x[9],a2_x[8],a2_x[7],a2_x[6],a2_x[5],a2_x[4],a2_x[3],a2_x[2],a2_x[1],a2_x[0]};
wire [1:0] a2addx = {a2addx_1,a2addx_0};
wire [23:0] address_ = {address[23],address[22],address[21],address[20],
address[19],address[18],address[17],address[16],address[15],address[14],address[13],address[12],address[11],address[10],
address[9],address[8],address[7],address[6],address[5],address[4],address[3],address[2],address[1],address[0]};
wire [7:0] dcomp = {dcomp_7,dcomp_6,dcomp_5,dcomp_4,dcomp_3,dcomp_2,dcomp_1,dcomp_0};
wire [31:0] gpu_din_ = {gpu_din[31],gpu_din[30],
gpu_din[29],gpu_din[28],gpu_din[27],gpu_din[26],gpu_din[25],gpu_din[24],gpu_din[23],gpu_din[22],gpu_din[21],gpu_din[20],
gpu_din[19],gpu_din[18],gpu_din[17],gpu_din[16],gpu_din[15],gpu_din[14],gpu_din[13],gpu_din[12],gpu_din[11],gpu_din[10],
gpu_din[9],gpu_din[8],gpu_din[7],gpu_din[6],gpu_din[5],gpu_din[4],gpu_din[3],gpu_din[2],gpu_din[1],gpu_din[0]};
wire [2:0] pixa = {pixa_2,pixa_1,pixa_0};
wire [7:0] srcd = {srcd_7,srcd_6,srcd_5,srcd_4,srcd_3,srcd_2,srcd_1,srcd_0};
wire [3:0] zcomp = {zcomp_3,zcomp_2,zcomp_1,zcomp_0};

_state state_inst
(
	.blit_addr_out /* BUS */ (blit_addr_out_[23:0]),
	.blit_addr_oe /* BUS */ (blit_addr_oe),
	.justify_out /* BUS */ (justify_out),
	.justify_oe /* BUS */ (justify_oe),
	.justify_in /* BUS */ (justify_in),
	.mreq_out /* BUS */ (mreq_out),
	.mreq_oe /* BUS */ (mreq_oe),
	.mreq_in /* BUS */ (mreq_in),
	.width_out /* BUS */ (width_out[3:0]),
	.width_oe /* BUS */ (width_0_oe),
	.read_out /* BUS */ (read_out),
	.read_oe /* BUS */ (read_oe),
	.read_in /* BUS */ (read_in),
	.gpu_dout_out /* BUS */ (gpu_dout_out[31:0]),
	.gpu_dout_oe /* BUS */ (gpu_dout_0_oe),
	.a1fracldi /* OUT */ (a1fracldi),
	.a1ptrldi /* OUT */ (a1ptrldi),
	.a2ptrldi /* OUT */ (a2ptrldi),
	.addasel /* OUT */ (addasel[2:0]),
	.addbsel /* OUT */ (addbsel[1:0]),
	.addqsel /* OUT */ (addqsel),
	.adda_xconst /* OUT */ (adda_xconst[2:0]),
	.adda_yconst /* OUT */ (adda_yconst),
	.addareg /* OUT */ (addareg),
	.apipe /* OUT */ (apipe),
	.blit_breq /* OUT */ (blit_breq[1:0]),
	.blit_int /* OUT */ (blit_int),
	.cmpdst /* OUT */ (cmpdst),
	.daddasel /* OUT */ (daddasel[2:0]),
	.daddbsel /* OUT */ (daddbsel[2:0]),
	.daddmode /* OUT */ (daddmode[2:0]),
	.data_ena /* OUT */ (data_ena),
	.data_sel /* OUT */ (data_sel[1:0]),
	.dbinh_n /* OUT */ (dbinh_n[7:0]),
	.dend /* OUT */ (dend[5:0]),
	.dpipe /* OUT */ (dpipe[1:0]),
	.dstart /* OUT */ (dstart[5:0]),
	.dstdread /* OUT */ (dstdread),
	.dstzread /* OUT */ (dstzread),
	.gena2 /* OUT */ (gena2),
	.lfu_func /* OUT */ (lfu_func[3:0]),
	.daddq_sel /* OUT */ (daddq_sel),
	.modx /* OUT */ (modx[2:0]),
	.patdadd /* OUT */ (patdadd),
	.patfadd /* OUT */ (patfadd),
	.phrase_mode /* OUT */ (phrase_mode),
	.reset_n /* OUT */ (reset_n),
	.srcdread /* OUT */ (srcdread),
	.srcshift /* OUT */ (srcshift[5:0]),
	.srcz1add /* OUT */ (srcz1add),
	.srcz2add /* OUT */ (srcz2add),
	.srczread /* OUT */ (srczread),
	.suba_x /* OUT */ (suba_x),
	.suba_y /* OUT */ (suba_y),
	.zaddr /* OUT */ (zaddr),
	.zmode /* OUT */ (zmode[2:0]),
	.zpipe /* OUT */ (zpipe[1:0]),
	.a1_outside /* IN */ (a1_outside),
	.a1_pixsize /* IN */ (a1_pixsize[2:0]),
	.a1_win_x /* IN */ (a1_win_x_[14:0]),
	.a1_x /* IN */ (a1_x_[15:0]),
	.a1addx /* IN */ (a1addx[1:0]),
	.a1addy /* IN */ (a1addy),
	.a1xsign /* IN */ (a1xsign),
	.a1ysign /* IN */ (a1ysign),
	.a2_pixsize /* IN */ (a2_pixsize[2:0]),
	.a2_x /* IN */ (a2_x_[15:0]),
	.a2addx /* IN */ (a2addx[1:0]),
	.a2addy /* IN */ (a2addy),
	.a2xsign /* IN */ (a2xsign),
	.a2ysign /* IN */ (a2ysign),
	.ack /* IN */ (ack),
	.address /* IN */ (address_[23:0]),
	.big_pix /* IN */ (big_pix),
	.blit_back /* IN */ (blit_back),
	.clk /* IN */ (clk),
	.cmdld /* IN */ (cmdld),
	.countld /* IN */ (countld),
	.dcomp /* IN */ (dcomp[7:0]),
	.gpu_din /* IN */ (gpu_din_[31:0]),
	.pixa /* IN */ (pixa[2:0]),
	.srcd /* IN */ (srcd[7:0]),
	.statrd /* IN */ (statrd),
	.stopld /* IN */ (stopld),
	.xreset_n /* IN */ (xreset_n),
	.zcomp /* IN */ (zcomp[3:0]),
	.sys_clk(sys_clk) // Generated
);

endmodule
