module sboard
(
	output [0:5] dsta,
	output sdatreq,
	output dstrwen_n,
	output [0:31] dstwd,
	output resaddrldi,
	output sbwait,
	output [0:5] srca,
	output srcaddrldi,
	output srcrwen_n,
	output [0:31] srcwd,
	input clk,
	input datack,
	input datwe,
	input datwe_raw,
	input del_xld,
	input div_activei,
	input div_instr,
	input div_start,
	input [0:5] dstanwi,
	input [0:5] dstat,
	input dstrrd,
	input dstrrdi,
	input dstrwr,
	input dstrwri,
	input dstwen,
	input exe,
	input flag_depend,
	input flagld,
	input gate_active,
	input [0:31] immdata,
	input immld,
	input immwri,
	input insexei,
	input [0:31] load_data,
	input [0:31] mem_data,
	input memrw,
	input mtx_dover,
	input precomp,
	input [0:31] quotient,
	input reset_n,
	input reswr,
	input [0:31] result,
	input [0:5] srcanwi,
	input [0:31] srcdp,
	input srcrrd,
	input xld_ready,
	input sys_clk // Generated
);
wire [5:0] dsta_;
assign {dsta[5],dsta[4],dsta[3],dsta[2],dsta[1],dsta[0]} = dsta_[5:0];
wire [31:0] dstwd_;
assign {dstwd[31],dstwd[30],
dstwd[29],dstwd[28],dstwd[27],dstwd[26],dstwd[25],dstwd[24],dstwd[23],dstwd[22],dstwd[21],dstwd[20],
dstwd[19],dstwd[18],dstwd[17],dstwd[16],dstwd[15],dstwd[14],dstwd[13],dstwd[12],dstwd[11],dstwd[10],
dstwd[9],dstwd[8],dstwd[7],dstwd[6],dstwd[5],dstwd[4],dstwd[3],dstwd[2],dstwd[1],dstwd[0]} = dstwd_[31:0];
wire [5:0] srca_;
assign {srca[5],srca[4],srca[3],srca[2],srca[1],srca[0]} = srca_[5:0];
wire [31:0] srcwd_;
assign {srcwd[31],srcwd[30],
srcwd[29],srcwd[28],srcwd[27],srcwd[26],srcwd[25],srcwd[24],srcwd[23],srcwd[22],srcwd[21],srcwd[20],
srcwd[19],srcwd[18],srcwd[17],srcwd[16],srcwd[15],srcwd[14],srcwd[13],srcwd[12],srcwd[11],srcwd[10],
srcwd[9],srcwd[8],srcwd[7],srcwd[6],srcwd[5],srcwd[4],srcwd[3],srcwd[2],srcwd[1],srcwd[0]} = srcwd_[31:0];
wire [5:0] dstanwi_ = {dstanwi[5],dstanwi[4],dstanwi[3],dstanwi[2],dstanwi[1],dstanwi[0]};
wire [5:0] dstat_ = {dstat[5],dstat[4],dstat[3],dstat[2],dstat[1],dstat[0]};
wire [31:0] immdata_ = {immdata[31],immdata[30],
immdata[29],immdata[28],immdata[27],immdata[26],immdata[25],immdata[24],immdata[23],immdata[22],immdata[21],immdata[20],
immdata[19],immdata[18],immdata[17],immdata[16],immdata[15],immdata[14],immdata[13],immdata[12],immdata[11],immdata[10],
immdata[9],immdata[8],immdata[7],immdata[6],immdata[5],immdata[4],immdata[3],immdata[2],immdata[1],immdata[0]};
wire [31:0] load_data_ = {load_data[31],load_data[30],
load_data[29],load_data[28],load_data[27],load_data[26],load_data[25],load_data[24],load_data[23],load_data[22],load_data[21],load_data[20],
load_data[19],load_data[18],load_data[17],load_data[16],load_data[15],load_data[14],load_data[13],load_data[12],load_data[11],load_data[10],
load_data[9],load_data[8],load_data[7],load_data[6],load_data[5],load_data[4],load_data[3],load_data[2],load_data[1],load_data[0]};
wire [31:0] mem_data_ = {mem_data[31],mem_data[30],
mem_data[29],mem_data[28],mem_data[27],mem_data[26],mem_data[25],mem_data[24],mem_data[23],mem_data[22],mem_data[21],mem_data[20],
mem_data[19],mem_data[18],mem_data[17],mem_data[16],mem_data[15],mem_data[14],mem_data[13],mem_data[12],mem_data[11],mem_data[10],
mem_data[9],mem_data[8],mem_data[7],mem_data[6],mem_data[5],mem_data[4],mem_data[3],mem_data[2],mem_data[1],mem_data[0]};
wire [31:0] quotient_ = {quotient[31],quotient[30],
quotient[29],quotient[28],quotient[27],quotient[26],quotient[25],quotient[24],quotient[23],quotient[22],quotient[21],quotient[20],
quotient[19],quotient[18],quotient[17],quotient[16],quotient[15],quotient[14],quotient[13],quotient[12],quotient[11],quotient[10],
quotient[9],quotient[8],quotient[7],quotient[6],quotient[5],quotient[4],quotient[3],quotient[2],quotient[1],quotient[0]};
wire [31:0] result_ = {result[31],result[30],
result[29],result[28],result[27],result[26],result[25],result[24],result[23],result[22],result[21],result[20],
result[19],result[18],result[17],result[16],result[15],result[14],result[13],result[12],result[11],result[10],
result[9],result[8],result[7],result[6],result[5],result[4],result[3],result[2],result[1],result[0]};
wire [5:0] srcanwi_ = {srcanwi[5],srcanwi[4],srcanwi[3],srcanwi[2],srcanwi[1],srcanwi[0]};
wire [31:0] srcdp_ = {srcdp[31],srcdp[30],
srcdp[29],srcdp[28],srcdp[27],srcdp[26],srcdp[25],srcdp[24],srcdp[23],srcdp[22],srcdp[21],srcdp[20],
srcdp[19],srcdp[18],srcdp[17],srcdp[16],srcdp[15],srcdp[14],srcdp[13],srcdp[12],srcdp[11],srcdp[10],
srcdp[9],srcdp[8],srcdp[7],srcdp[6],srcdp[5],srcdp[4],srcdp[3],srcdp[2],srcdp[1],srcdp[0]};
_sboard sboard_inst
(
	.dsta /* OUT */ (dsta_[5:0]),
	.sdatreq /* OUT */ (sdatreq),
	.dstrwen_n /* OUT */ (dstrwen_n),
	.dstwd /* OUT */ (dstwd_[31:0]),
	.resaddrldi /* OUT */ (resaddrldi),
	.sbwait /* OUT */ (sbwait),
	.srca /* OUT */ (srca_[5:0]),
	.srcaddrldi /* OUT */ (srcaddrldi),
	.srcrwen_n /* OUT */ (srcrwen_n),
	.srcwd /* OUT */ (srcwd_[31:0]),
	.clk /* IN */ (clk),
	.datack /* IN */ (datack),
	.datwe /* IN */ (datwe),
	.datwe_raw /* IN */ (datwe_raw),
	.del_xld /* IN */ (del_xld),
	.div_activei /* IN */ (div_activei),
	.div_instr /* IN */ (div_instr),
	.div_start /* IN */ (div_start),
	.dstanwi /* IN */ (dstanwi_[5:0]),
	.dstat /* IN */ (dstat_[5:0]),
	.dstrrd /* IN */ (dstrrd),
	.dstrrdi /* IN */ (dstrrdi),
	.dstrwr /* IN */ (dstrwr),
	.dstrwri /* IN */ (dstrwri),
	.dstwen /* IN */ (dstwen),
	.exe /* IN */ (exe),
	.flag_depend /* IN */ (flag_depend),
	.flagld /* IN */ (flagld),
	.gate_active /* IN */ (gate_active),
	.immdata /* IN */ (immdata_[31:0]),
	.immld /* IN */ (immld),
	.immwri /* IN */ (immwri),
	.insexei /* IN */ (insexei),
	.load_data /* IN */ (load_data_[31:0]),
	.mem_data /* IN */ (mem_data_[31:0]),
	.memrw /* IN */ (memrw),
	.mtx_dover /* IN */ (mtx_dover),
	.precomp /* IN */ (precomp),
	.quotient /* IN */ (quotient_[31:0]),
	.reset_n /* IN */ (reset_n),
	.reswr /* IN */ (reswr),
	.result /* IN */ (result_[31:0]),
	.srcanwi /* IN */ (srcanwi_[5:0]),
	.srcdp /* IN */ (srcdp_[31:0]),
	.srcrrd /* IN */ (srcrrd),
	.xld_ready /* IN */ (xld_ready),
	.sys_clk(sys_clk) // Generated
);
endmodule
