module ins_exec
(
	output [0:31] gpu_data_out,
	output [0:31] gpu_data_oe,
	input [0:31] gpu_data_in,
	output gpu_dout_3_out,
	output gpu_dout_3_oe,
	input gpu_dout_3_in,
	output gpu_dout_4_out,
	output gpu_dout_4_oe,
	input gpu_dout_4_in,
	output gpu_dout_5_out,
	output gpu_dout_5_oe,
	input gpu_dout_5_in,
	output gpu_dout_6_out,
	output gpu_dout_6_oe,
	input gpu_dout_6_in,
	output gpu_dout_7_out,
	output gpu_dout_7_oe,
	input gpu_dout_7_in,
	output gpu_dout_8_out,
	output gpu_dout_8_oe,
	input gpu_dout_8_in,
	output gpu_dout_9_out,
	output gpu_dout_9_oe,
	input gpu_dout_9_in,
	output gpu_dout_10_out,
	output gpu_dout_10_oe,
	input gpu_dout_10_in,
	output gpu_dout_11_out,
	output gpu_dout_11_oe,
	input gpu_dout_11_in,
	output gpu_dout_12_out,
	output gpu_dout_12_oe,
	input gpu_dout_12_in,
	output gpu_dout_13_out,
	output gpu_dout_13_oe,
	input gpu_dout_13_in,
	output gpu_dout_14_out,
	output gpu_dout_14_oe,
	input gpu_dout_14_in,
	output gpu_dout_16_out,
	output gpu_dout_16_oe,
	input gpu_dout_16_in,
	output gpu_dout_17_out,
	output gpu_dout_17_oe,
	input gpu_dout_17_in,
	output gpu_dout_18_out,
	output gpu_dout_18_oe,
	input gpu_dout_18_in,
	output gpu_dout_19_out,
	output gpu_dout_19_oe,
	input gpu_dout_19_in,
	output gpu_dout_20_out,
	output gpu_dout_20_oe,
	input gpu_dout_20_in,
	output gpu_dout_21_out,
	output gpu_dout_21_oe,
	input gpu_dout_21_in,
	output gpu_dout_22_out,
	output gpu_dout_22_oe,
	input gpu_dout_22_in,
	output gpu_dout_23_out,
	output gpu_dout_23_oe,
	input gpu_dout_23_in,
	output gpu_dout_24_out,
	output gpu_dout_24_oe,
	input gpu_dout_24_in,
	output gpu_dout_25_out,
	output gpu_dout_25_oe,
	input gpu_dout_25_in,
	output gpu_dout_26_out,
	output gpu_dout_26_oe,
	input gpu_dout_26_in,
	output gpu_dout_27_out,
	output gpu_dout_27_oe,
	input gpu_dout_27_in,
	output gpu_dout_28_out,
	output gpu_dout_28_oe,
	input gpu_dout_28_in,
	output gpu_dout_29_out,
	output gpu_dout_29_oe,
	input gpu_dout_29_in,
	output gpu_dout_30_out,
	output gpu_dout_30_oe,
	input gpu_dout_30_in,
	output gpu_dout_31_out,
	output gpu_dout_31_oe,
	input gpu_dout_31_in,
	output [0:2] alufunc,
	output brlmux_0,
	output brlmux_1,
	output [0:23] dataddr,
	output datreq,
	output datweb,
	output datwe_raw,
	output div_instr,
	output div_start,
	output [0:5] dstanwi,
	output [0:5] dstat,
	output dstdgate,
	output dstrrd,
	output dstrrdi,
	output dstrwr,
	output dstrwri,
	output dstwen,
	output exe,
	output flag_depend,
	output flagld,
	output [0:31] immdata,
	output immld,
	output immwri,
	output insexei,
	output locden,
	output [0:31] locsrc,
	output macop,
	output memrw,
	output msize_0,
	output msize_1,
	output mtx_dover,
	output multsel,
	output multsign,
	output pabort,
	output precomp,
	output [0:21] progaddr,
	output progreq,
	output resld,
	output ressel_0,
	output ressel_1,
	output ressel_2,
	output reswr,
	output rev_sub,
	output satsz_0,
	output satsz_1,
	output srcrrd,
	output single_stop,
	output [0:5] srcanwi,
	input big_instr,
	input carry_flag,
	input clk,
	input clkb,
	input tlw,
	input datack,
	input dbgrd,
	input div_activei,
	input external,
	input flagrd,
	input flagwr,
	input gate_active,
	input go,
	input [0:31] gpu_din,
	input gpu_irq_0,
	input gpu_irq_1,
	input gpu_irq_2,
	input gpu_irq_3,
	input gpu_irq_4,
	input gpu_irq_5, // jerry only
	input mtxawr,
	input mtxcwr,
	input nega_flag,
	input pcrd,
	input pcwr,
	input progack,
	input resaddrldi,
	input reset_n,
	input [0:31] result,
	input sbwait,
	input sdatreq,
	input single_go,
	input single_step,
	input srcaddrldi,
	input [0:31] srcd,
	input [0:31] srcdp,
	input [0:31] srcdpa,
	input statrd,
	input zero_flag,
	input sys_clk // Generated
);
parameter JERRY = 0;

wire [31:0] gpu_data_out_;
assign {gpu_data_out[31],gpu_data_out[30],
gpu_data_out[29],gpu_data_out[28],gpu_data_out[27],gpu_data_out[26],gpu_data_out[25],gpu_data_out[24],gpu_data_out[23],gpu_data_out[22],gpu_data_out[21],gpu_data_out[20],
gpu_data_out[19],gpu_data_out[18],gpu_data_out[17],gpu_data_out[16],gpu_data_out[15],gpu_data_out[14],gpu_data_out[13],gpu_data_out[12],gpu_data_out[11],gpu_data_out[10],
gpu_data_out[9],gpu_data_out[8],gpu_data_out[7],gpu_data_out[6],gpu_data_out[5],gpu_data_out[4],gpu_data_out[3],gpu_data_out[2],gpu_data_out[1],gpu_data_out[0]} = gpu_data_out_[31:0];
assign {gpu_data_oe[31],gpu_data_oe[30],
gpu_data_oe[29],gpu_data_oe[28],gpu_data_oe[27],gpu_data_oe[26],gpu_data_oe[25],gpu_data_oe[24],gpu_data_oe[23],gpu_data_oe[22],gpu_data_oe[21],gpu_data_oe[20],
gpu_data_oe[19],gpu_data_oe[18],gpu_data_oe[17],gpu_data_oe[16],gpu_data_oe[15],gpu_data_oe[14],gpu_data_oe[13],gpu_data_oe[12],gpu_data_oe[11],gpu_data_oe[10],
gpu_data_oe[9],gpu_data_oe[8],gpu_data_oe[7],gpu_data_oe[6],gpu_data_oe[5],gpu_data_oe[4],gpu_data_oe[3],gpu_data_oe[2],gpu_data_oe[1]} = {31{gpu_data_oe[0]}};
wire [31:0] gpu_data_in_ = {gpu_data_in[31],gpu_data_in[30],
gpu_data_in[29],gpu_data_in[28],gpu_data_in[27],gpu_data_in[26],gpu_data_in[25],gpu_data_in[24],gpu_data_in[23],gpu_data_in[22],gpu_data_in[21],gpu_data_in[20],
gpu_data_in[19],gpu_data_in[18],gpu_data_in[17],gpu_data_in[16],gpu_data_in[15],gpu_data_in[14],gpu_data_in[13],gpu_data_in[12],gpu_data_in[11],gpu_data_in[10],
gpu_data_in[9],gpu_data_in[8],gpu_data_in[7],gpu_data_in[6],gpu_data_in[5],gpu_data_in[4],gpu_data_in[3],gpu_data_in[2],gpu_data_in[1],gpu_data_in[0]};
wire [31:3] gpu_dout_out;
assign {gpu_dout_31_out,gpu_dout_30_out,
gpu_dout_29_out,gpu_dout_28_out,gpu_dout_27_out,gpu_dout_26_out,gpu_dout_25_out,gpu_dout_24_out,gpu_dout_23_out,gpu_dout_22_out,gpu_dout_21_out,gpu_dout_20_out,
gpu_dout_19_out,gpu_dout_18_out,gpu_dout_17_out,gpu_dout_16_out} = gpu_dout_out[31:16];
assign {gpu_dout_14_out,gpu_dout_13_out,gpu_dout_12_out,gpu_dout_11_out,gpu_dout_10_out,
gpu_dout_9_out,gpu_dout_8_out,gpu_dout_7_out,gpu_dout_6_out,gpu_dout_5_out,gpu_dout_4_out,gpu_dout_3_out} = gpu_dout_out[14:3];
assign {gpu_dout_31_oe,gpu_dout_30_oe,
gpu_dout_29_oe,gpu_dout_28_oe,gpu_dout_27_oe,gpu_dout_26_oe,gpu_dout_25_oe,gpu_dout_24_oe,gpu_dout_23_oe,gpu_dout_22_oe,gpu_dout_21_oe,gpu_dout_20_oe,
gpu_dout_19_oe,gpu_dout_18_oe,gpu_dout_17_oe} = {15{gpu_dout_16_oe}};
assign {gpu_dout_14_oe,gpu_dout_13_oe,gpu_dout_12_oe,gpu_dout_11_oe,gpu_dout_5_oe,gpu_dout_4_oe} = {6{gpu_dout_3_oe}};
assign {gpu_dout_10_oe,gpu_dout_9_oe,gpu_dout_8_oe,gpu_dout_7_oe} = {4{gpu_dout_6_oe}};

wire [2:0] alufunc_;
assign {alufunc[2],alufunc[1],alufunc[0]} = alufunc_[2:0];
wire [1:0] brlmux;
assign {brlmux_1,brlmux_0} = brlmux[1:0];
wire [23:0] dataddr_;
assign {dataddr[23],dataddr[22],dataddr[21],dataddr[20],
dataddr[19],dataddr[18],dataddr[17],dataddr[16],dataddr[15],dataddr[14],dataddr[13],dataddr[12],dataddr[11],dataddr[10],
dataddr[9],dataddr[8],dataddr[7],dataddr[6],dataddr[5],dataddr[4],dataddr[3],dataddr[2],dataddr[1],dataddr[0]} = dataddr_[23:0];
wire [5:0] dstanwi_;
assign {dstanwi[5],dstanwi[4],dstanwi[3],dstanwi[2],dstanwi[1],dstanwi[0]} = dstanwi_[5:0];
wire [5:0] dstat_;
assign {dstat[5],dstat[4],dstat[3],dstat[2],dstat[1],dstat[0]} = dstat_[5:0];
wire [31:0] immdata_;
assign {immdata[31],immdata[30],
immdata[29],immdata[28],immdata[27],immdata[26],immdata[25],immdata[24],immdata[23],immdata[22],immdata[21],immdata[20],
immdata[19],immdata[18],immdata[17],immdata[16],immdata[15],immdata[14],immdata[13],immdata[12],immdata[11],immdata[10],
immdata[9],immdata[8],immdata[7],immdata[6],immdata[5],immdata[4],immdata[3],immdata[2],immdata[1],immdata[0]} = immdata_[31:0];
wire [31:0] locsrc_;
assign {locsrc[31],locsrc[30],
locsrc[29],locsrc[28],locsrc[27],locsrc[26],locsrc[25],locsrc[24],locsrc[23],locsrc[22],locsrc[21],locsrc[20],
locsrc[19],locsrc[18],locsrc[17],locsrc[16],locsrc[15],locsrc[14],locsrc[13],locsrc[12],locsrc[11],locsrc[10],
locsrc[9],locsrc[8],locsrc[7],locsrc[6],locsrc[5],locsrc[4],locsrc[3],locsrc[2],locsrc[1],locsrc[0]} = locsrc_[31:0];
wire [1:0] msize;
assign {msize_1,msize_0} = msize[1:0];
wire [21:0] progaddr_;
assign {progaddr[21],progaddr[20],
progaddr[19],progaddr[18],progaddr[17],progaddr[16],progaddr[15],progaddr[14],progaddr[13],progaddr[12],progaddr[11],progaddr[10],
progaddr[9],progaddr[8],progaddr[7],progaddr[6],progaddr[5],progaddr[4],progaddr[3],progaddr[2],progaddr[1],progaddr[0]} = progaddr_[21:0];
wire [2:0] ressel;
assign {ressel_2,ressel_1,ressel_0} = ressel[2:0];
wire [1:0] satsz;
assign {satsz_1,satsz_0} = satsz[1:0];
wire [5:0] srcanwi_;
assign {srcanwi[5],srcanwi[4],srcanwi[3],srcanwi[2],srcanwi[1],srcanwi[0]} = srcanwi_[5:0];
wire [31:0] gpu_din_ = {gpu_din[31],gpu_din[30],
gpu_din[29],gpu_din[28],gpu_din[27],gpu_din[26],gpu_din[25],gpu_din[24],gpu_din[23],gpu_din[22],gpu_din[21],gpu_din[20],
gpu_din[19],gpu_din[18],gpu_din[17],gpu_din[16],gpu_din[15],gpu_din[14],gpu_din[13],gpu_din[12],gpu_din[11],gpu_din[10],
gpu_din[9],gpu_din[8],gpu_din[7],gpu_din[6],gpu_din[5],gpu_din[4],gpu_din[3],gpu_din[2],gpu_din[1],gpu_din[0]};
wire [5:0] gpu_irq = {gpu_irq_5,gpu_irq_4,gpu_irq_3,gpu_irq_2,gpu_irq_1,gpu_irq_0};
wire [31:0] result_ = {result[31],result[30],
result[29],result[28],result[27],result[26],result[25],result[24],result[23],result[22],result[21],result[20],
result[19],result[18],result[17],result[16],result[15],result[14],result[13],result[12],result[11],result[10],
result[9],result[8],result[7],result[6],result[5],result[4],result[3],result[2],result[1],result[0]};
wire [31:0] srcd_ = {srcd[31],srcd[30],
srcd[29],srcd[28],srcd[27],srcd[26],srcd[25],srcd[24],srcd[23],srcd[22],srcd[21],srcd[20],
srcd[19],srcd[18],srcd[17],srcd[16],srcd[15],srcd[14],srcd[13],srcd[12],srcd[11],srcd[10],
srcd[9],srcd[8],srcd[7],srcd[6],srcd[5],srcd[4],srcd[3],srcd[2],srcd[1],srcd[0]};
wire [31:0] srcdp_ = {srcdp[31],srcdp[30],
srcdp[29],srcdp[28],srcdp[27],srcdp[26],srcdp[25],srcdp[24],srcdp[23],srcdp[22],srcdp[21],srcdp[20],
srcdp[19],srcdp[18],srcdp[17],srcdp[16],srcdp[15],srcdp[14],srcdp[13],srcdp[12],srcdp[11],srcdp[10],
srcdp[9],srcdp[8],srcdp[7],srcdp[6],srcdp[5],srcdp[4],srcdp[3],srcdp[2],srcdp[1],srcdp[0]};
wire [31:0] srcdpa_ = {srcdpa[31],srcdpa[30],
srcdpa[29],srcdpa[28],srcdpa[27],srcdpa[26],srcdpa[25],srcdpa[24],srcdpa[23],srcdpa[22],srcdpa[21],srcdpa[20],
srcdpa[19],srcdpa[18],srcdpa[17],srcdpa[16],srcdpa[15],srcdpa[14],srcdpa[13],srcdpa[12],srcdpa[11],srcdpa[10],
srcdpa[9],srcdpa[8],srcdpa[7],srcdpa[6],srcdpa[5],srcdpa[4],srcdpa[3],srcdpa[2],srcdpa[1],srcdpa[0]};
_ins_exec #(.JERRY(JERRY)) ins_exec_inst
(
	.gpu_data_out /* BUS */ (gpu_data_out_[31:0]),
	.gpu_data_oe /* BUS */ (gpu_data_oe[0]),
	.gpu_data_in /* BUS */ (gpu_data_in_[31:0]),
	.gpu_dout_out /* BUS */ (gpu_dout_out[31:3]), //15 not used
	.gpu_dout_14_3_oe /* BUS */ (gpu_dout_3_oe),
	.gpu_dout_10_6_oe /* BUS */ (gpu_dout_6_oe),
	.gpu_dout_31_16_oe /* BUS */ (gpu_dout_16_oe),
	.alufunc /* OUT */ (alufunc_[2:0]),
	.brlmux /* OUT */ (brlmux[1:0]),
	.dataddr /* OUT */ (dataddr_[23:0]),
	.datreq /* OUT */ (datreq),
	.datweb /* OUT */ (datweb),
	.datwe_raw /* OUT */ (datwe_raw),
	.div_instr /* OUT */ (div_instr),
	.div_start /* OUT */ (div_start),
	.dstanwi /* OUT */ (dstanwi_[5:0]),
	.dstat /* OUT */ (dstat_[5:0]),
	.dstdgate /* OUT */ (dstdgate),
	.dstrrd /* OUT */ (dstrrd),
	.dstrrdi /* OUT */ (dstrrdi),
	.dstrwr /* OUT */ (dstrwr),
	.dstrwri /* OUT */ (dstrwri),
	.dstwen /* OUT */ (dstwen),
	.exe /* OUT */ (exe),
	.flag_depend /* OUT */ (flag_depend),
	.flagld /* OUT */ (flagld),
	.immdata /* OUT */ (immdata_[31:0]),
	.immld /* OUT */ (immld),
	.immwri /* OUT */ (immwri),
	.insexei /* OUT */ (insexei),
	.locden /* OUT */ (locden),
	.locsrc /* OUT */ (locsrc_[31:0]),
	.macop /* OUT */ (macop),
	.memrw /* OUT */ (memrw),
	.msize /* OUT */ (msize[1:0]),
	.mtx_dover /* OUT */ (mtx_dover),
	.multsel /* OUT */ (multsel),
	.multsign /* OUT */ (multsign),
	.pabort /* OUT */ (pabort),
	.precomp /* OUT */ (precomp),
	.progaddr /* OUT */ (progaddr_[21:0]),
	.progreq /* OUT */ (progreq),
	.resld /* OUT */ (resld),
	.ressel /* OUT */ (ressel[2:0]),
	.reswr /* OUT */ (reswr),
	.rev_sub /* OUT */ (rev_sub),
	.satsz /* OUT */ (satsz[1:0]),
	.srcrrd /* OUT */ (srcrrd),
	.single_stop /* OUT */ (single_stop),
	.srcanwi /* OUT */ (srcanwi_[5:0]),
	.big_instr /* IN */ (big_instr),
	.carry_flag /* IN */ (carry_flag),
	.clk /* IN */ (clk),
	.clkb /* IN */ (clkb),
	.tlw /* IN */ (tlw),
	.datack /* IN */ (datack),
	.dbgrd /* IN */ (dbgrd),
	.div_activei /* IN */ (div_activei),
	.external /* IN */ (external),
	.flagrd /* IN */ (flagrd),
	.flagwr /* IN */ (flagwr),
	.gate_active /* IN */ (gate_active),
	.go /* IN */ (go),
	.gpu_din /* IN */ (gpu_din_[31:0]),
	.gpu_irq /* IN */ (gpu_irq[5:0]),
	.mtxawr /* IN */ (mtxawr),
	.mtxcwr /* IN */ (mtxcwr),
	.nega_flag /* IN */ (nega_flag),
	.pcrd /* IN */ (pcrd),
	.pcwr /* IN */ (pcwr),
	.progack /* IN */ (progack),
	.resaddrldi /* IN */ (resaddrldi),
	.reset_n /* IN */ (reset_n),
	.result /* IN */ (result_[31:0]),
	.sbwait /* IN */ (sbwait),
	.sdatreq /* IN */ (sdatreq),
	.single_go /* IN */ (single_go),
	.single_step /* IN */ (single_step),
	.srcaddrldi /* IN */ (srcaddrldi),
	.srcd /* IN */ (srcd_[31:0]),
	.srcdp /* IN */ (srcdp_[31:0]),
	.srcdpa /* IN */ (srcdpa_[31:0]),
	.statrd /* IN */ (statrd),
	.zero_flag /* IN */ (zero_flag),
	.sys_clk(sys_clk) // Generated
);

endmodule
