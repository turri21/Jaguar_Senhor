/* verilator lint_off LITENDIAN */
//`include "defs.v"

module j_dsp
(
	input ima_0,
	input ima_1,
	input ima_2,
	input ima_3,
	input ima_4,
	input ima_5,
	input ima_6,
	input ima_7,
	input ima_8,
	input ima_9,
	input ima_10,
	input ima_11,
	input ima_12,
	input ima_13,
	input ima_14,
	input ima_15,
	input dout_0,
	input dout_1,
	input dout_2,
	input dout_3,
	input dout_4,
	input dout_5,
	input dout_6,
	input dout_7,
	input dout_8,
	input dout_9,
	input dout_10,
	input dout_11,
	input dout_12,
	input dout_13,
	input dout_14,
	input dout_15,
	input dout_16,
	input dout_17,
	input dout_18,
	input dout_19,
	input dout_20,
	input dout_21,
	input dout_22,
	input dout_23,
	input dout_24,
	input dout_25,
	input dout_26,
	input dout_27,
	input dout_28,
	input dout_29,
	input dout_30,
	input dout_31,
	input tlw_a,
	input tlw_b,
	input tlw_c,
	input ack,
	input gpu_back,
	input reset_n,
	input clk,
	input eint_n_0,
	input eint_n_1,
	input tint_0,
	input tint_1,
	input i2int,
	input iord,
	input iowr,
	input tlw,
	output gpu_breq,
	output dma_breq,
	output cpu_int,
	output wdata_0,
	output wdata_1,
	output wdata_2,
	output wdata_3,
	output wdata_4,
	output wdata_5,
	output wdata_6,
	output wdata_7,
	output wdata_8,
	output wdata_9,
	output wdata_10,
	output wdata_11,
	output wdata_12,
	output wdata_13,
	output wdata_14,
	output wdata_15,
	output wdata_16,
	output wdata_17,
	output wdata_18,
	output wdata_19,
	output wdata_20,
	output wdata_21,
	output wdata_22,
	output wdata_23,
	output wdata_24,
	output wdata_25,
	output wdata_26,
	output wdata_27,
	output wdata_28,
	output wdata_29,
	output wdata_30,
	output wdata_31,
	output a_0,
	output a_1,
	output a_2,
	output a_3,
	output a_4,
	output a_5,
	output a_6,
	output a_7,
	output a_8,
	output a_9,
	output a_10,
	output a_11,
	output a_12,
	output a_13,
	output a_14,
	output a_15,
	output a_16,
	output a_17,
	output a_18,
	output a_19,
	output a_20,
	output a_21,
	output a_22,
	output a_23,
	output width_0,
	output width_1,
	output width_2,
	output read,
	output mreq,
	output dacw_0,
	output dacw_1,
	output gpu_din_0,
	output gpu_din_1,
	output gpu_din_2,
	output gpu_din_3,
	output gpu_din_4,
	output gpu_din_5,
	output gpu_din_6,
	output gpu_din_7,
	output gpu_din_8,
	output gpu_din_9,
	output gpu_din_10,
	output gpu_din_11,
	output gpu_din_12,
	output gpu_din_13,
	output gpu_din_14,
	output gpu_din_15,
	output i2sw_0,
	output i2sw_1,
	output i2sw_2,
	output i2sw_3,
	output i2sr_0,
	output i2sr_1,
	output i2sr_2,
	output dr_0_out,
	output dr_0_oe,
	input dr_0_in,
	output dr_1_out,
	output dr_1_oe,
	input dr_1_in,
	output dr_2_out,
	output dr_2_oe,
	input dr_2_in,
	output dr_3_out,
	output dr_3_oe,
	input dr_3_in,
	output dr_4_out,
	output dr_4_oe,
	input dr_4_in,
	output dr_5_out,
	output dr_5_oe,
	input dr_5_in,
	output dr_6_out,
	output dr_6_oe,
	input dr_6_in,
	output dr_7_out,
	output dr_7_oe,
	input dr_7_in,
	output dr_8_out,
	output dr_8_oe,
	input dr_8_in,
	output dr_9_out,
	output dr_9_oe,
	input dr_9_in,
	output dr_10_out,
	output dr_10_oe,
	input dr_10_in,
	output dr_11_out,
	output dr_11_oe,
	input dr_11_in,
	output dr_12_out,
	output dr_12_oe,
	input dr_12_in,
	output dr_13_out,
	output dr_13_oe,
	input dr_13_in,
	output dr_14_out,
	output dr_14_oe,
	input dr_14_in,
	output dr_15_out,
	output dr_15_oe,
	input dr_15_in,
	output gpu_dout_o_0_out,
	output gpu_dout_o_0_oe,
	input gpu_dout_o_0_in,
	output gpu_dout_o_1_out,
	output gpu_dout_o_1_oe,
	input gpu_dout_o_1_in,
	output gpu_dout_o_2_out,
	output gpu_dout_o_2_oe,
	input gpu_dout_o_2_in,
	output gpu_dout_o_3_out,
	output gpu_dout_o_3_oe,
	input gpu_dout_o_3_in,
	output gpu_dout_o_4_out,
	output gpu_dout_o_4_oe,
	input gpu_dout_o_4_in,
	output gpu_dout_o_5_out,
	output gpu_dout_o_5_oe,
	input gpu_dout_o_5_in,
	output gpu_dout_o_6_out,
	output gpu_dout_o_6_oe,
	input gpu_dout_o_6_in,
	output gpu_dout_o_7_out,
	output gpu_dout_o_7_oe,
	input gpu_dout_o_7_in,
	output gpu_dout_o_8_out,
	output gpu_dout_o_8_oe,
	input gpu_dout_o_8_in,
	output gpu_dout_o_9_out,
	output gpu_dout_o_9_oe,
	input gpu_dout_o_9_in,
	output gpu_dout_o_10_out,
	output gpu_dout_o_10_oe,
	input gpu_dout_o_10_in,
	output gpu_dout_o_11_out,
	output gpu_dout_o_11_oe,
	input gpu_dout_o_11_in,
	output gpu_dout_o_12_out,
	output gpu_dout_o_12_oe,
	input gpu_dout_o_12_in,
	output gpu_dout_o_13_out,
	output gpu_dout_o_13_oe,
	input gpu_dout_o_13_in,
	output gpu_dout_o_14_out,
	output gpu_dout_o_14_oe,
	input gpu_dout_o_14_in,
	output gpu_dout_o_15_out,
	output gpu_dout_o_15_oe,
	input gpu_dout_o_15_in,
	input sys_clk // Generated
);
wire [15:0] ima = {ima_15,ima_14,ima_13,ima_12,ima_11,ima_10,
ima_9,ima_8,ima_7,ima_6,ima_5,ima_4,ima_3,ima_2,ima_1,ima_0};
wire [31:0] dout = {dout_31,dout_30,
dout_29,dout_28,dout_27,dout_26,dout_25,dout_24,dout_23,dout_22,dout_21,dout_20,
dout_19,dout_18,dout_17,dout_16,dout_15,dout_14,dout_13,dout_12,dout_11,dout_10,
dout_9,dout_8,dout_7,dout_6,dout_5,dout_4,dout_3,dout_2,dout_1,dout_0};
wire [1:0] eint_n = {eint_n_1,eint_n_0};
wire [1:0] tint = {tint_1,tint_0};
wire [31:0] wdata;
assign {wdata_31,wdata_30,
wdata_29,wdata_28,wdata_27,wdata_26,wdata_25,wdata_24,wdata_23,wdata_22,wdata_21,wdata_20,
wdata_19,wdata_18,wdata_17,wdata_16,wdata_15,wdata_14,wdata_13,wdata_12,wdata_11,wdata_10,
wdata_9,wdata_8,wdata_7,wdata_6,wdata_5,wdata_4,wdata_3,wdata_2,wdata_1,wdata_0} = wdata[31:0];
wire [23:0] a;
assign {a_23,a_22,a_21,a_20,
a_19,a_18,a_17,a_16,a_15,a_14,a_13,a_12,a_11,a_10,
a_9,a_8,a_7,a_6,a_5,a_4,a_3,a_2,a_1,a_0} = a[23:0];
wire [2:0] width;
assign {width_2,width_1,width_0} = width[2:0];
wire [1:0] dacw;
assign {dacw_1,dacw_0} = dacw[1:0];
wire [15:0] gpu_din;
assign {gpu_din_15,gpu_din_14,gpu_din_13,gpu_din_12,gpu_din_11,gpu_din_10,
gpu_din_9,gpu_din_8,gpu_din_7,gpu_din_6,gpu_din_5,gpu_din_4,gpu_din_3,gpu_din_2,gpu_din_1,gpu_din_0} = gpu_din[15:0];
wire [15:0] dr_out;
assign {dr_15_out,dr_14_out,dr_13_out,dr_12_out,dr_11_out,dr_10_out,
dr_9_out,dr_8_out,dr_7_out,dr_6_out,dr_5_out,dr_4_out,dr_3_out,dr_2_out,dr_1_out,dr_0_out} = dr_out[15:0];
assign {dr_15_oe,dr_14_oe,dr_13_oe,dr_12_oe,dr_11_oe,dr_10_oe,
dr_9_oe,dr_8_oe,dr_7_oe,dr_6_oe,dr_5_oe,dr_4_oe,dr_3_oe,dr_2_oe,dr_1_oe} = {15{dr_0_oe}};
wire [15:0] gpu_dout_o_out;
assign {gpu_dout_o_15_out,gpu_dout_o_14_out,gpu_dout_o_13_out,gpu_dout_o_12_out,gpu_dout_o_11_out,gpu_dout_o_10_out,
gpu_dout_o_9_out,gpu_dout_o_8_out,gpu_dout_o_7_out,gpu_dout_o_6_out,gpu_dout_o_5_out,gpu_dout_o_4_out,gpu_dout_o_3_out,gpu_dout_o_2_out,gpu_dout_o_1_out,gpu_dout_o_0_out} = gpu_dout_o_out[15:0];
assign {gpu_dout_o_15_oe,gpu_dout_o_14_oe,gpu_dout_o_13_oe,gpu_dout_o_12_oe,gpu_dout_o_11_oe,gpu_dout_o_10_oe,
gpu_dout_o_9_oe,gpu_dout_o_8_oe,gpu_dout_o_7_oe,gpu_dout_o_6_oe,gpu_dout_o_5_oe,gpu_dout_o_4_oe,gpu_dout_o_3_oe,gpu_dout_o_2_oe,gpu_dout_o_1_oe} = {15{gpu_dout_o_0_oe}};
wire [15:0] gpu_dout_o_in = {gpu_dout_o_15_in,gpu_dout_o_14_in,gpu_dout_o_13_in,gpu_dout_o_12_in,gpu_dout_o_11_in,gpu_dout_o_10_in,
gpu_dout_o_9_in,gpu_dout_o_8_in,gpu_dout_o_7_in,gpu_dout_o_6_in,gpu_dout_o_5_in,gpu_dout_o_4_in,gpu_dout_o_3_in,gpu_dout_o_2_in,gpu_dout_o_1_in,gpu_dout_o_0_in};
_j_dsp dsp_inst
(
	.ima /* IN */ (ima[15:0]),		// I/O address.
	.dout /* IN */ (dout[31:0]),		// slave write / master read data.
	.ack /* IN */ (ack),					// co-processor memory acknowledge.
	.gpu_back /* IN */ (gpu_back),			// GPU normal bus acknowledge.
	.reset_n /* IN */ (reset_n),		// system reset.
	.clk /* IN */ (clk),					// system clock.
	.eint_n /* IN */ (eint_n[1:0]),		// external interrupts.
	.tint /* IN */ (tint[1:0]),			// timer interrupts.
	.i2int /* IN */ (i2int),			// I2S interrupt.
	.iord /* IN */ (iord),			// Look-ahead I/O read strobe for GPU.
	.iowr /* IN */ (iowr),			// Look-ahead I/O write strobe for GPU.
	.tlw /* IN */ (tlw),					// Transparent latch write enable timing.
	.tlw_a        (tlw_a),
	.tlw_b        (tlw_b),
	.tlw_c        (tlw_c),
	.gpu_breq /* OUT */ (gpu_breq),	// GPU normal bus request.
	.dma_breq /* OUT */ (dma_breq),	// GPU high-priority bus request.
	.cpu_int /* OUT */ (cpu_int),			// GPU interrupt to CPU.
	.wdata /* OUT */ (wdata[31:0]),			// master write data bus.
	.a /* OUT */ (a[23:0]),				// master cycle address bus.
	.width /* OUT */ (width[2:0]),			// master cycle cycle width (in bytes).
	.read /* OUT */ (read),				// master cycle read request.
	.mreq /* OUT */ (mreq),				// master cycle request.
	.dacw /* OUT */ (dacw[1:0]),			// internal DAC write strobes.
	.gpu_din /* OUT */ (gpu_din[15:0]),	// internal I/O write data.
	.i2sw_0 /* OUT */ (i2sw_0),    // LTXD Left transmit data F1A148 WO.
	.i2sw_1 /* OUT */ (i2sw_1),    // RTXD Right transmit data F1A14C WO.
	.i2sw_2 /* OUT */ (i2sw_2),    // SCLK Serial Clock Frequency F1A150 WO.
	.i2sw_3 /* OUT */ (i2sw_3),    // SMODE Serial Mode F1A154 WO.
	.i2sr_0 /* OUT */ (i2sr_0),		// internal I2S read strobes.
	.i2sr_1 /* OUT */ (i2sr_1),
	.i2sr_2 /* OUT */ (i2sr_2),
	.dr_out /* BUS */ (dr_out[15:0]),	// I/O read data (busses split, and OE added, for Verilog translation).
	.dr_oe /* BUS */ (dr_0_oe),
	.gpu_dout_o_out /* BUS */ (gpu_dout_o_out[15:0]),	// read data from internal peripherals (GE - renamed).
	.gpu_dout_o_oe /* BUS */ (gpu_dout_o_0_oe),
	.gpu_dout_o_in /* BUS */ (gpu_dout_o_in[15:0]),
	.sys_clk(sys_clk) // Generated
);
endmodule
