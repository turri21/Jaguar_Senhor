module gpu_ctrl
(
	output gpu_dout_0_out,
	output gpu_dout_0_oe,
	input gpu_dout_0_in,
	output gpu_dout_1_out,
	output gpu_dout_1_oe,
	input gpu_dout_1_in,
	output gpu_dout_2_out,
	output gpu_dout_2_oe,
	input gpu_dout_2_in,
	output gpu_dout_3_out,
	output gpu_dout_3_oe,
	input gpu_dout_3_in,
	output gpu_dout_4_out,
	output gpu_dout_4_oe,
	input gpu_dout_4_in,
	output gpu_dout_5_out,
	output gpu_dout_5_oe,
	input gpu_dout_5_in,
	output gpu_dout_11_out,
	output gpu_dout_11_oe,
	input gpu_dout_11_in,
	output gpu_dout_12_out,
	output gpu_dout_12_oe,
	input gpu_dout_12_in,
	output gpu_dout_13_out,
	output gpu_dout_13_oe,
	input gpu_dout_13_in,
	output gpu_dout_14_out,
	output gpu_dout_14_oe,
	input gpu_dout_14_in,
	output gpu_dout_15_out,
	output gpu_dout_15_oe,
	input gpu_dout_15_in,
	output bus_hog,
	output cpu_int,
	output go,
	output gpu_irq_0,
	output single_go,
	output single_step,
	input clk,
	input ctrlwr,
	input ctrlwrgo,
	input [0:31] gpu_din,
	input reset_n,
	input single_stop,
	input statrd,
	input sys_clk // Generated
);
wire [15:0] gpu_dout_out;
assign {gpu_dout_15_out,gpu_dout_14_out,gpu_dout_13_out,gpu_dout_12_out,gpu_dout_11_out} = gpu_dout_out[15:11];
assign {gpu_dout_5_out,gpu_dout_4_out,gpu_dout_3_out,gpu_dout_2_out,gpu_dout_1_out,gpu_dout_0_out} = gpu_dout_out[5:0];
assign {gpu_dout_15_oe,gpu_dout_14_oe,gpu_dout_13_oe,gpu_dout_12_oe} = {4{gpu_dout_11_oe}};
assign {gpu_dout_5_oe,gpu_dout_4_oe,gpu_dout_3_oe,gpu_dout_2_oe,gpu_dout_1_oe} = {5{gpu_dout_0_oe}};
wire [31:0] gpu_din_ = {gpu_din[31],gpu_din[30],
gpu_din[29],gpu_din[28],gpu_din[27],gpu_din[26],gpu_din[25],gpu_din[24],gpu_din[23],gpu_din[22],gpu_din[21],gpu_din[20],
gpu_din[19],gpu_din[18],gpu_din[17],gpu_din[16],gpu_din[15],gpu_din[14],gpu_din[13],gpu_din[12],gpu_din[11],gpu_din[10],
gpu_din[9],gpu_din[8],gpu_din[7],gpu_din[6],gpu_din[5],gpu_din[4],gpu_din[3],gpu_din[2],gpu_din[1],gpu_din[0]};
_gpu_ctrl gpu_ctrl_inst
(
	.gpu_dout_out /* BUS */ (gpu_dout_out[15:0]),
	.gpu_dout_5_0_oe /* BUS */ (gpu_dout_0_oe), 
	.gpu_dout_15_11_oe /* BUS */ (gpu_dout_11_oe),
	.bus_hog /* OUT */ (bus_hog),
	.cpu_int /* OUT */ (cpu_int),
	.go /* OUT */ (go),
	.gpu_irq_0 /* OUT */ (gpu_irq_0),
	.single_go /* OUT */ (single_go),
	.single_step /* OUT */ (single_step),
	.clk /* IN */ (clk),
	.ctrlwr /* IN */ (ctrlwr),
	.ctrlwrgo /* IN */ (ctrlwrgo),
	.gpu_din /* IN */ (gpu_din_[31:0]),
	.reset_n /* IN */ (reset_n),
	.single_stop /* IN */ (single_stop),
	.statrd /* IN */ (statrd),
	.sys_clk(sys_clk) // Generated
);
endmodule
