//`include "defs.v"
// altera message_off 10036

module wbk
(
	input d_14,
	input d_15,
	input d_16,
	input d_17,
	input d_18,
	input d_19,
	input d_20,
	input d_21,
	input d_22,
	input d_23,
	input d_43,
	input d_44,
	input d_45,
	input d_46,
	input d_47,
	input d_48,
	input d_49,
	input d_50,
	input d_51,
	input d_52,
	input d_53,
	input d_54,
	input d_55,
	input d_56,
	input d_57,
	input d_58,
	input d_59,
	input d_60,
	input d_61,
	input d_62,
	input d_63,
	input obld_0,
	input obld_2,
	input dwidth_0,
	input dwidth_1,
	input dwidth_2,
	input dwidth_3,
	input dwidth_4,
	input dwidth_5,
	input dwidth_6,
	input dwidth_7,
	input dwidth_8,
	input dwidth_9,
	input vscale_0,
	input vscale_1,
	input vscale_2,
	input vscale_3,
	input vscale_4,
	input vscale_5,
	input vscale_6,
	input vscale_7,
	input clk,
	input resetl,
	input scaled,
	input wbkstart,
	output newdata_0,
	output newdata_1,
	output newdata_2,
	output newdata_3,
	output newdata_4,
	output newdata_5,
	output newdata_6,
	output newdata_7,
	output newdata_8,
	output newdata_9,
	output newdata_10,
	output newdata_11,
	output newdata_12,
	output newdata_13,
	output newdata_14,
	output newdata_15,
	output newdata_16,
	output newdata_17,
	output newdata_18,
	output newdata_19,
	output newdata_20,
	output newheight_0,
	output newheight_1,
	output newheight_2,
	output newheight_3,
	output newheight_4,
	output newheight_5,
	output newheight_6,
	output newheight_7,
	output newheight_8,
	output newheight_9,
	output newrem_0,
	output newrem_1,
	output newrem_2,
	output newrem_3,
	output newrem_4,
	output newrem_5,
	output newrem_6,
	output newrem_7,
	output heightnz,
	output wbkdone,
	input sys_clk // Generated
);
wire [63:0] d = {d_63,d_62,d_61,d_60,
d_59,d_58,d_57,d_56,d_55,d_54,d_53,d_52,d_51,d_50,
d_49,d_48,d_47,d_46,d_45,d_44,d_43,
19'h0,
d_23,d_22,d_21,d_20,
d_19,d_18,d_17,d_16,d_15,d_14,
14'h0};
wire [7:0] vscale = {vscale_7,vscale_6,vscale_5,vscale_4,vscale_3,vscale_2,vscale_1,vscale_0};
wire [9:0] dwidth = {dwidth_9,dwidth_8,dwidth_7,dwidth_6,dwidth_5,dwidth_4,dwidth_3,dwidth_2,dwidth_1,dwidth_0};
wire [20:0] newdata;
assign {newdata_20,
newdata_19,newdata_18,newdata_17,newdata_16,newdata_15,newdata_14,newdata_13,newdata_12,newdata_11,newdata_10,
newdata_9,newdata_8,newdata_7,newdata_6,newdata_5,newdata_4,newdata_3,newdata_2,newdata_1,newdata_0} = newdata[20:0];
wire [9:0] newheight;
assign {newheight_9,newheight_8,newheight_7,newheight_6,newheight_5,newheight_4,newheight_3,newheight_2,newheight_1,newheight_0} = newheight[9:0];
wire [7:0] newrem;
assign {newrem_7,newrem_6,newrem_5,newrem_4,newrem_3,newrem_2,newrem_1,newrem_0} = newrem[7:0];
_wbk wbk_inst
(
	.d /* IN */ (d[63:0]),// only d[23:14] and d[63:43] used
	.obld_0 /* IN */ (obld_0),
	.obld_2 /* IN */ (obld_2),
	.dwidth /* IN */ (dwidth[9:0]),
	.vscale /* IN */ (vscale[7:0]),
	.clk /* IN */ (clk),
	.resetl /* IN */ (resetl),
	.scaled /* IN */ (scaled),
	.wbkstart /* IN */ (wbkstart),
	.newdata /* OUT */ (newdata[20:0]),
	.newheight /* OUT */ (newheight[9:0]),
	.newrem /* OUT */ (newrem[7:0]),
	.heightnz /* OUT */ (heightnz),
	.wbkdone /* OUT */ (wbkdone),
	.sys_clk(sys_clk) // Generated
);
endmodule
