module graphics
(
	input ima_0,
	input ima_1,
	input ima_2,
	input ima_3,
	input ima_4,
	input ima_5,
	input ima_6,
	input ima_7,
	input ima_8,
	input ima_9,
	input ima_10,
	input ima_11,
	input ima_12,
	input ima_13,
	input ima_14,
	input ima_15,
	input dwrite_0,
	input dwrite_1,
	input dwrite_2,
	input dwrite_3,
	input dwrite_4,
	input dwrite_5,
	input dwrite_6,
	input dwrite_7,
	input dwrite_8,
	input dwrite_9,
	input dwrite_10,
	input dwrite_11,
	input dwrite_12,
	input dwrite_13,
	input dwrite_14,
	input dwrite_15,
	input dwrite_16,
	input dwrite_17,
	input dwrite_18,
	input dwrite_19,
	input dwrite_20,
	input dwrite_21,
	input dwrite_22,
	input dwrite_23,
	input dwrite_24,
	input dwrite_25,
	input dwrite_26,
	input dwrite_27,
	input dwrite_28,
	input dwrite_29,
	input dwrite_30,
	input dwrite_31,
	input ack,
	input blit_back,
	input gpu_back,
	input reset_n,
	input clk,
	input tlw,
	input dint,
	input gpu_irq_3,
	input gpu_irq_2,
	input iord,
	input iowr,
	input reset_lock,
	input data_0,
	input data_1,
	input data_2,
	input data_3,
	input data_4,
	input data_5,
	input data_6,
	input data_7,
	input data_8,
	input data_9,
	input data_10,
	input data_11,
	input data_12,
	input data_13,
	input data_14,
	input data_15,
	input data_16,
	input data_17,
	input data_18,
	input data_19,
	input data_20,
	input data_21,
	input data_22,
	input data_23,
	input data_24,
	input data_25,
	input data_26,
	input data_27,
	input data_28,
	input data_29,
	input data_30,
	input data_31,
	input data_32,
	input data_33,
	input data_34,
	input data_35,
	input data_36,
	input data_37,
	input data_38,
	input data_39,
	input data_40,
	input data_41,
	input data_42,
	input data_43,
	input data_44,
	input data_45,
	input data_46,
	input data_47,
	input data_48,
	input data_49,
	input data_50,
	input data_51,
	input data_52,
	input data_53,
	input data_54,
	input data_55,
	input data_56,
	input data_57,
	input data_58,
	input data_59,
	input data_60,
	input data_61,
	input data_62,
	input data_63,
	input at_1,
	output blit_breq_0,
	output blit_breq_1,
	output gpu_breq,
	output dma_breq,
	output cpu_int,
	output lock,
	output wdata_0_out,
	output wdata_0_oe,
	input wdata_0_in,
	output wdata_1_out,
	output wdata_1_oe,
	input wdata_1_in,
	output wdata_2_out,
	output wdata_2_oe,
	input wdata_2_in,
	output wdata_3_out,
	output wdata_3_oe,
	input wdata_3_in,
	output wdata_4_out,
	output wdata_4_oe,
	input wdata_4_in,
	output wdata_5_out,
	output wdata_5_oe,
	input wdata_5_in,
	output wdata_6_out,
	output wdata_6_oe,
	input wdata_6_in,
	output wdata_7_out,
	output wdata_7_oe,
	input wdata_7_in,
	output wdata_8_out,
	output wdata_8_oe,
	input wdata_8_in,
	output wdata_9_out,
	output wdata_9_oe,
	input wdata_9_in,
	output wdata_10_out,
	output wdata_10_oe,
	input wdata_10_in,
	output wdata_11_out,
	output wdata_11_oe,
	input wdata_11_in,
	output wdata_12_out,
	output wdata_12_oe,
	input wdata_12_in,
	output wdata_13_out,
	output wdata_13_oe,
	input wdata_13_in,
	output wdata_14_out,
	output wdata_14_oe,
	input wdata_14_in,
	output wdata_15_out,
	output wdata_15_oe,
	input wdata_15_in,
	output wdata_16_out,
	output wdata_16_oe,
	input wdata_16_in,
	output wdata_17_out,
	output wdata_17_oe,
	input wdata_17_in,
	output wdata_18_out,
	output wdata_18_oe,
	input wdata_18_in,
	output wdata_19_out,
	output wdata_19_oe,
	input wdata_19_in,
	output wdata_20_out,
	output wdata_20_oe,
	input wdata_20_in,
	output wdata_21_out,
	output wdata_21_oe,
	input wdata_21_in,
	output wdata_22_out,
	output wdata_22_oe,
	input wdata_22_in,
	output wdata_23_out,
	output wdata_23_oe,
	input wdata_23_in,
	output wdata_24_out,
	output wdata_24_oe,
	input wdata_24_in,
	output wdata_25_out,
	output wdata_25_oe,
	input wdata_25_in,
	output wdata_26_out,
	output wdata_26_oe,
	input wdata_26_in,
	output wdata_27_out,
	output wdata_27_oe,
	input wdata_27_in,
	output wdata_28_out,
	output wdata_28_oe,
	input wdata_28_in,
	output wdata_29_out,
	output wdata_29_oe,
	input wdata_29_in,
	output wdata_30_out,
	output wdata_30_oe,
	input wdata_30_in,
	output wdata_31_out,
	output wdata_31_oe,
	input wdata_31_in,
	output wdata_32_out,
	output wdata_32_oe,
	input wdata_32_in,
	output wdata_33_out,
	output wdata_33_oe,
	input wdata_33_in,
	output wdata_34_out,
	output wdata_34_oe,
	input wdata_34_in,
	output wdata_35_out,
	output wdata_35_oe,
	input wdata_35_in,
	output wdata_36_out,
	output wdata_36_oe,
	input wdata_36_in,
	output wdata_37_out,
	output wdata_37_oe,
	input wdata_37_in,
	output wdata_38_out,
	output wdata_38_oe,
	input wdata_38_in,
	output wdata_39_out,
	output wdata_39_oe,
	input wdata_39_in,
	output wdata_40_out,
	output wdata_40_oe,
	input wdata_40_in,
	output wdata_41_out,
	output wdata_41_oe,
	input wdata_41_in,
	output wdata_42_out,
	output wdata_42_oe,
	input wdata_42_in,
	output wdata_43_out,
	output wdata_43_oe,
	input wdata_43_in,
	output wdata_44_out,
	output wdata_44_oe,
	input wdata_44_in,
	output wdata_45_out,
	output wdata_45_oe,
	input wdata_45_in,
	output wdata_46_out,
	output wdata_46_oe,
	input wdata_46_in,
	output wdata_47_out,
	output wdata_47_oe,
	input wdata_47_in,
	output wdata_48_out,
	output wdata_48_oe,
	input wdata_48_in,
	output wdata_49_out,
	output wdata_49_oe,
	input wdata_49_in,
	output wdata_50_out,
	output wdata_50_oe,
	input wdata_50_in,
	output wdata_51_out,
	output wdata_51_oe,
	input wdata_51_in,
	output wdata_52_out,
	output wdata_52_oe,
	input wdata_52_in,
	output wdata_53_out,
	output wdata_53_oe,
	input wdata_53_in,
	output wdata_54_out,
	output wdata_54_oe,
	input wdata_54_in,
	output wdata_55_out,
	output wdata_55_oe,
	input wdata_55_in,
	output wdata_56_out,
	output wdata_56_oe,
	input wdata_56_in,
	output wdata_57_out,
	output wdata_57_oe,
	input wdata_57_in,
	output wdata_58_out,
	output wdata_58_oe,
	input wdata_58_in,
	output wdata_59_out,
	output wdata_59_oe,
	input wdata_59_in,
	output wdata_60_out,
	output wdata_60_oe,
	input wdata_60_in,
	output wdata_61_out,
	output wdata_61_oe,
	input wdata_61_in,
	output wdata_62_out,
	output wdata_62_oe,
	input wdata_62_in,
	output wdata_63_out,
	output wdata_63_oe,
	input wdata_63_in,
	output a_0_out,
	output a_0_oe,
	input a_0_in,
	output a_1_out,
	output a_1_oe,
	input a_1_in,
	output a_2_out,
	output a_2_oe,
	input a_2_in,
	output a_3_out,
	output a_3_oe,
	input a_3_in,
	output a_4_out,
	output a_4_oe,
	input a_4_in,
	output a_5_out,
	output a_5_oe,
	input a_5_in,
	output a_6_out,
	output a_6_oe,
	input a_6_in,
	output a_7_out,
	output a_7_oe,
	input a_7_in,
	output a_8_out,
	output a_8_oe,
	input a_8_in,
	output a_9_out,
	output a_9_oe,
	input a_9_in,
	output a_10_out,
	output a_10_oe,
	input a_10_in,
	output a_11_out,
	output a_11_oe,
	input a_11_in,
	output a_12_out,
	output a_12_oe,
	input a_12_in,
	output a_13_out,
	output a_13_oe,
	input a_13_in,
	output a_14_out,
	output a_14_oe,
	input a_14_in,
	output a_15_out,
	output a_15_oe,
	input a_15_in,
	output a_16_out,
	output a_16_oe,
	input a_16_in,
	output a_17_out,
	output a_17_oe,
	input a_17_in,
	output a_18_out,
	output a_18_oe,
	input a_18_in,
	output a_19_out,
	output a_19_oe,
	input a_19_in,
	output a_20_out,
	output a_20_oe,
	input a_20_in,
	output a_21_out,
	output a_21_oe,
	input a_21_in,
	output a_22_out,
	output a_22_oe,
	input a_22_in,
	output a_23_out,
	output a_23_oe,
	input a_23_in,
	output width_0_out,
	output width_0_oe,
	input width_0_in,
	output width_1_out,
	output width_1_oe,
	input width_1_in,
	output width_2_out,
	output width_2_oe,
	input width_2_in,
	output width_3_out,
	output width_3_oe,
	input width_3_in,
	output read_out,
	output read_oe,
	input read_in,
	output mreq_out,
	output mreq_oe,
	input mreq_in,
	output dr_0_out,
	output dr_0_oe,
	input dr_0_in,
	output dr_1_out,
	output dr_1_oe,
	input dr_1_in,
	output dr_2_out,
	output dr_2_oe,
	input dr_2_in,
	output dr_3_out,
	output dr_3_oe,
	input dr_3_in,
	output dr_4_out,
	output dr_4_oe,
	input dr_4_in,
	output dr_5_out,
	output dr_5_oe,
	input dr_5_in,
	output dr_6_out,
	output dr_6_oe,
	input dr_6_in,
	output dr_7_out,
	output dr_7_oe,
	input dr_7_in,
	output dr_8_out,
	output dr_8_oe,
	input dr_8_in,
	output dr_9_out,
	output dr_9_oe,
	input dr_9_in,
	output dr_10_out,
	output dr_10_oe,
	input dr_10_in,
	output dr_11_out,
	output dr_11_oe,
	input dr_11_in,
	output dr_12_out,
	output dr_12_oe,
	input dr_12_in,
	output dr_13_out,
	output dr_13_oe,
	input dr_13_in,
	output dr_14_out,
	output dr_14_oe,
	input dr_14_in,
	output dr_15_out,
	output dr_15_oe,
	input dr_15_in,
	output justify_out,
	output justify_oe,
	input justify_in,
	input sys_clk // Generated
);
wire [15:0] ima = {ima_15,ima_14,ima_13,ima_12,ima_11,ima_10,
ima_9,ima_8,ima_7,ima_6,ima_5,ima_4,ima_3,ima_2,ima_1,ima_0};
wire [31:0] dwrite = {dwrite_31,dwrite_30,
dwrite_29,dwrite_28,dwrite_27,dwrite_26,dwrite_25,dwrite_24,dwrite_23,dwrite_22,dwrite_21,dwrite_20,
dwrite_19,dwrite_18,dwrite_17,dwrite_16,dwrite_15,dwrite_14,dwrite_13,dwrite_12,dwrite_11,dwrite_10,
dwrite_9,dwrite_8,dwrite_7,dwrite_6,dwrite_5,dwrite_4,dwrite_3,dwrite_2,dwrite_1,dwrite_0};
wire [3:2] gpu_irq = {gpu_irq_3,gpu_irq_2};//3 2
wire [63:0] data = {data_63,data_62,data_61,data_60,
data_59,data_58,data_57,data_56,data_55,data_54,data_53,data_52,data_51,data_50,
data_49,data_48,data_47,data_46,data_45,data_44,data_43,data_42,data_41,data_40,
data_39,data_38,data_37,data_36,data_35,data_34,data_33,data_32,data_31,data_30,
data_29,data_28,data_27,data_26,data_25,data_24,data_23,data_22,data_21,data_20,
data_19,data_18,data_17,data_16,data_15,data_14,data_13,data_12,data_11,data_10,
data_9,data_8,data_7,data_6,data_5,data_4,data_3,data_2,data_1,data_0};
wire [1:0] blit_breq;
assign {blit_breq_1,blit_breq_0} = blit_breq[1:0];
wire [63:0] wdata_out;
assign {wdata_63_out,wdata_62_out,wdata_61_out,wdata_60_out,
wdata_59_out,wdata_58_out,wdata_57_out,wdata_56_out,wdata_55_out,wdata_54_out,wdata_53_out,wdata_52_out,wdata_51_out,wdata_50_out,
wdata_49_out,wdata_48_out,wdata_47_out,wdata_46_out,wdata_45_out,wdata_44_out,wdata_43_out,wdata_42_out,wdata_41_out,wdata_40_out,
wdata_39_out,wdata_38_out,wdata_37_out,wdata_36_out,wdata_35_out,wdata_34_out,wdata_33_out,wdata_32_out,wdata_31_out,wdata_30_out,
wdata_29_out,wdata_28_out,wdata_27_out,wdata_26_out,wdata_25_out,wdata_24_out,wdata_23_out,wdata_22_out,wdata_21_out,wdata_20_out,
wdata_19_out,wdata_18_out,wdata_17_out,wdata_16_out,wdata_15_out,wdata_14_out,wdata_13_out,wdata_12_out,wdata_11_out,wdata_10_out,
wdata_9_out,wdata_8_out,wdata_7_out,wdata_6_out,wdata_5_out,wdata_4_out,wdata_3_out,wdata_2_out,wdata_1_out,wdata_0_out} = wdata_out[63:0];
assign {wdata_63_oe,wdata_62_oe,wdata_61_oe,wdata_60_oe,
wdata_59_oe,wdata_58_oe,wdata_57_oe,wdata_56_oe,wdata_55_oe,wdata_54_oe,wdata_53_oe,wdata_52_oe,wdata_51_oe,wdata_50_oe,
wdata_49_oe,wdata_48_oe,wdata_47_oe,wdata_46_oe,wdata_45_oe,wdata_44_oe,wdata_43_oe,wdata_42_oe,wdata_41_oe,wdata_40_oe,
wdata_39_oe,wdata_38_oe,wdata_37_oe,wdata_36_oe,wdata_35_oe,wdata_34_oe,wdata_33_oe} = {31{wdata_32_oe}};
assign {wdata_31_oe,wdata_30_oe,
wdata_29_oe,wdata_28_oe,wdata_27_oe,wdata_26_oe,wdata_25_oe,wdata_24_oe,wdata_23_oe,wdata_22_oe,wdata_21_oe,wdata_20_oe,
wdata_19_oe,wdata_18_oe,wdata_17_oe,wdata_16_oe,wdata_15_oe,wdata_14_oe,wdata_13_oe,wdata_12_oe,wdata_11_oe,wdata_10_oe,
wdata_9_oe,wdata_8_oe,wdata_7_oe,wdata_6_oe,wdata_5_oe,wdata_4_oe,wdata_3_oe,wdata_2_oe,wdata_1_oe} = {31{wdata_0_oe}};
wire [23:0] a_out;
assign {a_23_out,a_22_out,a_21_out,a_20_out,
a_19_out,a_18_out,a_17_out,a_16_out,a_15_out,a_14_out,a_13_out,a_12_out,a_11_out,a_10_out,
a_9_out,a_8_out,a_7_out,a_6_out,a_5_out,a_4_out,a_3_out,a_2_out,a_1_out,a_0_out} = a_out[23:0];
assign {a_23_oe,a_22_oe,a_21_oe,a_20_oe,
a_19_oe,a_18_oe,a_17_oe,a_16_oe,a_15_oe,a_14_oe,a_13_oe,a_12_oe,a_11_oe,a_10_oe,
a_9_oe,a_8_oe,a_7_oe,a_6_oe,a_5_oe,a_4_oe,a_3_oe,a_2_oe,a_1_oe} = {23{a_0_oe}};
wire [3:0] width_out;
assign {width_3_out,width_2_out,width_1_out,width_0_out} = width_out[3:0];
assign {width_3_oe,width_2_oe,width_1_oe} = {3{width_0_oe}};
wire [15:0] dr_out;
assign {dr_15_out,dr_14_out,dr_13_out,dr_12_out,dr_11_out,dr_10_out,
dr_9_out,dr_8_out,dr_7_out,dr_6_out,dr_5_out,dr_4_out,dr_3_out,dr_2_out,dr_1_out,dr_0_out} = dr_out[15:0];
assign {dr_15_oe,dr_14_oe,dr_13_oe,dr_12_oe,dr_11_oe,dr_10_oe,
dr_9_oe,dr_8_oe,dr_7_oe,dr_6_oe,dr_5_oe,dr_4_oe,dr_3_oe,dr_2_oe,dr_1_oe} = {15{dr_0_oe}};
_graphics gpu_inst
(
	.ima /* IN */ (ima[15:0]),
	.dwrite /* IN */ (dwrite[31:0]),
	.ack /* IN */ (ack),
	.blit_back /* IN */ (blit_back),
	.gpu_back /* IN */ (gpu_back),
	.reset_n /* IN */ (reset_n),
	.clk /* IN */ (clk),
	.tlw /* IN */ (tlw),
	.dint /* IN */ (dint),
	.gpu_irq /* IN */ (gpu_irq[3:2]),//3 2
	.iord /* IN */ (iord),
	.iowr /* IN */ (iowr),
	.reset_lock /* IN */ (reset_lock),
	.data /* IN */ (data[63:0]),
	.at_1 /* IN */ (at_1),
	.blit_breq /* OUT */ (blit_breq[1:0]),
	.gpu_breq /* OUT */ (gpu_breq),
	.dma_breq /* OUT */ (dma_breq),
	.cpu_int /* OUT */ (cpu_int),
	.lock /* OUT */ (lock),
	.wdata_out /* BUS */ (wdata_out[63:0]),
	.wdata_31_0_oe /* BUS */ (wdata_0_oe),
	.wdata_63_32_oe /* BUS */ (wdata_32_oe),
	.a_out /* BUS */ (a_out[23:0]),
	.a_oe /* BUS */ (a_0_oe),
	.a_15_in /* BUS */ (a_15_in),
	.width_out /* BUS */ (width_out[3:0]),
	.width_oe /* BUS */ (width_0_oe),
	.read_out /* BUS */ (read_out),
	.read_oe /* BUS */ (read_oe),
	.read_in /* BUS */ (read_in),
	.mreq_out /* BUS */ (mreq_out),
	.mreq_oe /* BUS */ (mreq_oe),
	.mreq_in /* BUS */ (mreq_in),
	.dr_out /* BUS */ (dr_out[15:0]),
	.dr_oe /* BUS */ (dr_0_oe),
	.justify_out /* BUS */ (justify_out),
	.justify_oe /* BUS */ (justify_oe),
	.justify_in /* BUS */ (justify_in),
	.sys_clk(sys_clk) // Generated
);

endmodule
