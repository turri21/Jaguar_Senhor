//`include "defs.v"

module osc4c
(
	output	z0,
	output	z1,
	input 	a
);

// I don't know what it does
assign z0 = a;
assign z1 = a;

endmodule
