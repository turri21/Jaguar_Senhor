module __data_mux
(
	output wdata_0_out,
	output wdata_0_oe,
	input wdata_0_in,
	output wdata_1_out,
	output wdata_1_oe,
	input wdata_1_in,
	output wdata_2_out,
	output wdata_2_oe,
	input wdata_2_in,
	output wdata_3_out,
	output wdata_3_oe,
	input wdata_3_in,
	output wdata_4_out,
	output wdata_4_oe,
	input wdata_4_in,
	output wdata_5_out,
	output wdata_5_oe,
	input wdata_5_in,
	output wdata_6_out,
	output wdata_6_oe,
	input wdata_6_in,
	output wdata_7_out,
	output wdata_7_oe,
	input wdata_7_in,
	output wdata_8_out,
	output wdata_8_oe,
	input wdata_8_in,
	output wdata_9_out,
	output wdata_9_oe,
	input wdata_9_in,
	output wdata_10_out,
	output wdata_10_oe,
	input wdata_10_in,
	output wdata_11_out,
	output wdata_11_oe,
	input wdata_11_in,
	output wdata_12_out,
	output wdata_12_oe,
	input wdata_12_in,
	output wdata_13_out,
	output wdata_13_oe,
	input wdata_13_in,
	output wdata_14_out,
	output wdata_14_oe,
	input wdata_14_in,
	output wdata_15_out,
	output wdata_15_oe,
	input wdata_15_in,
	output wdata_16_out,
	output wdata_16_oe,
	input wdata_16_in,
	output wdata_17_out,
	output wdata_17_oe,
	input wdata_17_in,
	output wdata_18_out,
	output wdata_18_oe,
	input wdata_18_in,
	output wdata_19_out,
	output wdata_19_oe,
	input wdata_19_in,
	output wdata_20_out,
	output wdata_20_oe,
	input wdata_20_in,
	output wdata_21_out,
	output wdata_21_oe,
	input wdata_21_in,
	output wdata_22_out,
	output wdata_22_oe,
	input wdata_22_in,
	output wdata_23_out,
	output wdata_23_oe,
	input wdata_23_in,
	output wdata_24_out,
	output wdata_24_oe,
	input wdata_24_in,
	output wdata_25_out,
	output wdata_25_oe,
	input wdata_25_in,
	output wdata_26_out,
	output wdata_26_oe,
	input wdata_26_in,
	output wdata_27_out,
	output wdata_27_oe,
	input wdata_27_in,
	output wdata_28_out,
	output wdata_28_oe,
	input wdata_28_in,
	output wdata_29_out,
	output wdata_29_oe,
	input wdata_29_in,
	output wdata_30_out,
	output wdata_30_oe,
	input wdata_30_in,
	output wdata_31_out,
	output wdata_31_oe,
	input wdata_31_in,
	output wdata_32_out,
	output wdata_32_oe,
	input wdata_32_in,
	output wdata_33_out,
	output wdata_33_oe,
	input wdata_33_in,
	output wdata_34_out,
	output wdata_34_oe,
	input wdata_34_in,
	output wdata_35_out,
	output wdata_35_oe,
	input wdata_35_in,
	output wdata_36_out,
	output wdata_36_oe,
	input wdata_36_in,
	output wdata_37_out,
	output wdata_37_oe,
	input wdata_37_in,
	output wdata_38_out,
	output wdata_38_oe,
	input wdata_38_in,
	output wdata_39_out,
	output wdata_39_oe,
	input wdata_39_in,
	output wdata_40_out,
	output wdata_40_oe,
	input wdata_40_in,
	output wdata_41_out,
	output wdata_41_oe,
	input wdata_41_in,
	output wdata_42_out,
	output wdata_42_oe,
	input wdata_42_in,
	output wdata_43_out,
	output wdata_43_oe,
	input wdata_43_in,
	output wdata_44_out,
	output wdata_44_oe,
	input wdata_44_in,
	output wdata_45_out,
	output wdata_45_oe,
	input wdata_45_in,
	output wdata_46_out,
	output wdata_46_oe,
	input wdata_46_in,
	output wdata_47_out,
	output wdata_47_oe,
	input wdata_47_in,
	output wdata_48_out,
	output wdata_48_oe,
	input wdata_48_in,
	output wdata_49_out,
	output wdata_49_oe,
	input wdata_49_in,
	output wdata_50_out,
	output wdata_50_oe,
	input wdata_50_in,
	output wdata_51_out,
	output wdata_51_oe,
	input wdata_51_in,
	output wdata_52_out,
	output wdata_52_oe,
	input wdata_52_in,
	output wdata_53_out,
	output wdata_53_oe,
	input wdata_53_in,
	output wdata_54_out,
	output wdata_54_oe,
	input wdata_54_in,
	output wdata_55_out,
	output wdata_55_oe,
	input wdata_55_in,
	output wdata_56_out,
	output wdata_56_oe,
	input wdata_56_in,
	output wdata_57_out,
	output wdata_57_oe,
	input wdata_57_in,
	output wdata_58_out,
	output wdata_58_oe,
	input wdata_58_in,
	output wdata_59_out,
	output wdata_59_oe,
	input wdata_59_in,
	output wdata_60_out,
	output wdata_60_oe,
	input wdata_60_in,
	output wdata_61_out,
	output wdata_61_oe,
	input wdata_61_in,
	output wdata_62_out,
	output wdata_62_oe,
	input wdata_62_in,
	output wdata_63_out,
	output wdata_63_oe,
	input wdata_63_in,
	input [0:15] addq_0,
	input [0:15] addq_1,
	input [0:15] addq_2,
	input [0:15] addq_3,
	input big_pix,
	input [0:31] dstdlo,
	input [0:31] dstdhi,
	input [0:31] dstzlo,
	input [0:31] dstzhi,
	input data_sel_0,
	input data_sel_1,
	input data_ena,
	input dstart_0,
	input dstart_1,
	input dstart_2,
	input dstart_3,
	input dstart_4,
	input dstart_5,
	input dend_0,
	input dend_1,
	input dend_2,
	input dend_3,
	input dend_4,
	input dend_5,
	input dbinh_n_0,
	input dbinh_n_1,
	input dbinh_n_2,
	input dbinh_n_3,
	input dbinh_n_4,
	input dbinh_n_5,
	input dbinh_n_6,
	input dbinh_n_7,
	input [0:31] lfu_0,
	input [0:31] lfu_1,
	input [0:31] patd_0,
	input [0:31] patd_1,
	input phrase_mode,
	input [0:31] srczlo,
	input [0:31] srczhi
);
wire [63:0] wdata_out;
assign {wdata_63_out,wdata_62_out,wdata_61_out,wdata_60_out,
wdata_59_out,wdata_58_out,wdata_57_out,wdata_56_out,wdata_55_out,wdata_54_out,wdata_53_out,wdata_52_out,wdata_51_out,wdata_50_out,
wdata_49_out,wdata_48_out,wdata_47_out,wdata_46_out,wdata_45_out,wdata_44_out,wdata_43_out,wdata_42_out,wdata_41_out,wdata_40_out,
wdata_39_out,wdata_38_out,wdata_37_out,wdata_36_out,wdata_35_out,wdata_34_out,wdata_33_out,wdata_32_out,wdata_31_out,wdata_30_out,
wdata_29_out,wdata_28_out,wdata_27_out,wdata_26_out,wdata_25_out,wdata_24_out,wdata_23_out,wdata_22_out,wdata_21_out,wdata_20_out,
wdata_19_out,wdata_18_out,wdata_17_out,wdata_16_out,wdata_15_out,wdata_14_out,wdata_13_out,wdata_12_out,wdata_11_out,wdata_10_out,
wdata_9_out,wdata_8_out,wdata_7_out,wdata_6_out,wdata_5_out,wdata_4_out,wdata_3_out,wdata_2_out,wdata_1_out,wdata_0_out} = wdata_out[63:0];
assign {wdata_63_oe,wdata_62_oe,wdata_61_oe,wdata_60_oe,
wdata_59_oe,wdata_58_oe,wdata_57_oe,wdata_56_oe,wdata_55_oe,wdata_54_oe,wdata_53_oe,wdata_52_oe,wdata_51_oe,wdata_50_oe,
wdata_49_oe,wdata_48_oe,wdata_47_oe,wdata_46_oe,wdata_45_oe,wdata_44_oe,wdata_43_oe,wdata_42_oe,wdata_41_oe,wdata_40_oe,
wdata_39_oe,wdata_38_oe,wdata_37_oe,wdata_36_oe,wdata_35_oe,wdata_34_oe,wdata_33_oe,wdata_32_oe,wdata_31_oe,wdata_30_oe,
wdata_29_oe,wdata_28_oe,wdata_27_oe,wdata_26_oe,wdata_25_oe,wdata_24_oe,wdata_23_oe,wdata_22_oe,wdata_21_oe,wdata_20_oe,
wdata_19_oe,wdata_18_oe,wdata_17_oe,wdata_16_oe,wdata_15_oe,wdata_14_oe,wdata_13_oe,wdata_12_oe,wdata_11_oe,wdata_10_oe,
wdata_9_oe,wdata_8_oe,wdata_7_oe,wdata_6_oe,wdata_5_oe,wdata_4_oe,wdata_3_oe,wdata_2_oe,wdata_1_oe} = {63{wdata_0_oe}};
wire [15:0] addq_0_ = {addq_0[15],addq_0[14],addq_0[13],addq_0[12],addq_0[11],addq_0[10],
addq_0[9],addq_0[8],addq_0[7],addq_0[6],addq_0[5],addq_0[4],addq_0[3],addq_0[2],addq_0[1],addq_0[0]};
wire [15:0] addq_1_ = {addq_1[15],addq_1[14],addq_1[13],addq_1[12],addq_1[11],addq_1[10],
addq_1[9],addq_1[8],addq_1[7],addq_1[6],addq_1[5],addq_1[4],addq_1[3],addq_1[2],addq_1[1],addq_1[0]};
wire [15:0] addq_2_ = {addq_2[15],addq_2[14],addq_2[13],addq_2[12],addq_2[11],addq_2[10],
addq_2[9],addq_2[8],addq_2[7],addq_2[6],addq_2[5],addq_2[4],addq_2[3],addq_2[2],addq_2[1],addq_2[0]};
wire [15:0] addq_3_ = {addq_3[15],addq_3[14],addq_3[13],addq_3[12],addq_3[11],addq_3[10],
addq_3[9],addq_3[8],addq_3[7],addq_3[6],addq_3[5],addq_3[4],addq_3[3],addq_3[2],addq_3[1],addq_3[0]};
wire [31:0] dstdlo_ = {dstdlo[31],dstdlo[30],
dstdlo[29],dstdlo[28],dstdlo[27],dstdlo[26],dstdlo[25],dstdlo[24],dstdlo[23],dstdlo[22],dstdlo[21],dstdlo[20],
dstdlo[19],dstdlo[18],dstdlo[17],dstdlo[16],dstdlo[15],dstdlo[14],dstdlo[13],dstdlo[12],dstdlo[11],dstdlo[10],
dstdlo[9],dstdlo[8],dstdlo[7],dstdlo[6],dstdlo[5],dstdlo[4],dstdlo[3],dstdlo[2],dstdlo[1],dstdlo[0]};
wire [31:0] dstdhi_ = {dstdhi[31],dstdhi[30],
dstdhi[29],dstdhi[28],dstdhi[27],dstdhi[26],dstdhi[25],dstdhi[24],dstdhi[23],dstdhi[22],dstdhi[21],dstdhi[20],
dstdhi[19],dstdhi[18],dstdhi[17],dstdhi[16],dstdhi[15],dstdhi[14],dstdhi[13],dstdhi[12],dstdhi[11],dstdhi[10],
dstdhi[9],dstdhi[8],dstdhi[7],dstdhi[6],dstdhi[5],dstdhi[4],dstdhi[3],dstdhi[2],dstdhi[1],dstdhi[0]};
wire [31:0] dstzlo_ = {dstzlo[31],dstzlo[30],
dstzlo[29],dstzlo[28],dstzlo[27],dstzlo[26],dstzlo[25],dstzlo[24],dstzlo[23],dstzlo[22],dstzlo[21],dstzlo[20],
dstzlo[19],dstzlo[18],dstzlo[17],dstzlo[16],dstzlo[15],dstzlo[14],dstzlo[13],dstzlo[12],dstzlo[11],dstzlo[10],
dstzlo[9],dstzlo[8],dstzlo[7],dstzlo[6],dstzlo[5],dstzlo[4],dstzlo[3],dstzlo[2],dstzlo[1],dstzlo[0]};
wire [31:0] dstzhi_ = {dstzhi[31],dstzhi[30],
dstzhi[29],dstzhi[28],dstzhi[27],dstzhi[26],dstzhi[25],dstzhi[24],dstzhi[23],dstzhi[22],dstzhi[21],dstzhi[20],
dstzhi[19],dstzhi[18],dstzhi[17],dstzhi[16],dstzhi[15],dstzhi[14],dstzhi[13],dstzhi[12],dstzhi[11],dstzhi[10],
dstzhi[9],dstzhi[8],dstzhi[7],dstzhi[6],dstzhi[5],dstzhi[4],dstzhi[3],dstzhi[2],dstzhi[1],dstzhi[0]};
wire [1:0] data_sel = {data_sel_1,data_sel_0};
wire [5:0] dstart = {dstart_5,dstart_4,dstart_3,dstart_2,dstart_1,dstart_0};
wire [5:0] dend = {dend_5,dend_4,dend_3,dend_2,dend_1,dend_0};
wire [7:0] dbinh_n = {dbinh_n_7,dbinh_n_6,dbinh_n_5,dbinh_n_4,dbinh_n_3,dbinh_n_2,dbinh_n_1,dbinh_n_0};
wire [31:0] lfu_0_ = {lfu_0[31],lfu_0[30],
lfu_0[29],lfu_0[28],lfu_0[27],lfu_0[26],lfu_0[25],lfu_0[24],lfu_0[23],lfu_0[22],lfu_0[21],lfu_0[20],
lfu_0[19],lfu_0[18],lfu_0[17],lfu_0[16],lfu_0[15],lfu_0[14],lfu_0[13],lfu_0[12],lfu_0[11],lfu_0[10],
lfu_0[9],lfu_0[8],lfu_0[7],lfu_0[6],lfu_0[5],lfu_0[4],lfu_0[3],lfu_0[2],lfu_0[1],lfu_0[0]};
wire [31:0] lfu_1_ = {lfu_1[31],lfu_1[30],
lfu_1[29],lfu_1[28],lfu_1[27],lfu_1[26],lfu_1[25],lfu_1[24],lfu_1[23],lfu_1[22],lfu_1[21],lfu_1[20],
lfu_1[19],lfu_1[18],lfu_1[17],lfu_1[16],lfu_1[15],lfu_1[14],lfu_1[13],lfu_1[12],lfu_1[11],lfu_1[10],
lfu_1[9],lfu_1[8],lfu_1[7],lfu_1[6],lfu_1[5],lfu_1[4],lfu_1[3],lfu_1[2],lfu_1[1],lfu_1[0]};
wire [31:0] patd_0_ = {patd_0[31],patd_0[30],
patd_0[29],patd_0[28],patd_0[27],patd_0[26],patd_0[25],patd_0[24],patd_0[23],patd_0[22],patd_0[21],patd_0[20],
patd_0[19],patd_0[18],patd_0[17],patd_0[16],patd_0[15],patd_0[14],patd_0[13],patd_0[12],patd_0[11],patd_0[10],
patd_0[9],patd_0[8],patd_0[7],patd_0[6],patd_0[5],patd_0[4],patd_0[3],patd_0[2],patd_0[1],patd_0[0]};
wire [31:0] patd_1_ = {patd_1[31],patd_1[30],
patd_1[29],patd_1[28],patd_1[27],patd_1[26],patd_1[25],patd_1[24],patd_1[23],patd_1[22],patd_1[21],patd_1[20],
patd_1[19],patd_1[18],patd_1[17],patd_1[16],patd_1[15],patd_1[14],patd_1[13],patd_1[12],patd_1[11],patd_1[10],
patd_1[9],patd_1[8],patd_1[7],patd_1[6],patd_1[5],patd_1[4],patd_1[3],patd_1[2],patd_1[1],patd_1[0]};
wire [31:0] srczlo_ = {srczlo[31],srczlo[30],
srczlo[29],srczlo[28],srczlo[27],srczlo[26],srczlo[25],srczlo[24],srczlo[23],srczlo[22],srczlo[21],srczlo[20],
srczlo[19],srczlo[18],srczlo[17],srczlo[16],srczlo[15],srczlo[14],srczlo[13],srczlo[12],srczlo[11],srczlo[10],
srczlo[9],srczlo[8],srczlo[7],srczlo[6],srczlo[5],srczlo[4],srczlo[3],srczlo[2],srczlo[1],srczlo[0]};
wire [31:0] srczhi_ = {srczhi[31],srczhi[30],
srczhi[29],srczhi[28],srczhi[27],srczhi[26],srczhi[25],srczhi[24],srczhi[23],srczhi[22],srczhi[21],srczhi[20],
srczhi[19],srczhi[18],srczhi[17],srczhi[16],srczhi[15],srczhi[14],srczhi[13],srczhi[12],srczhi[11],srczhi[10],
srczhi[9],srczhi[8],srczhi[7],srczhi[6],srczhi[5],srczhi[4],srczhi[3],srczhi[2],srczhi[1],srczhi[0]};
_data_mux data_out_inst
(
	.wdata_out /* BUS */ (wdata_out[63:0]),
	.wdata_oe /* BUS */ (wdata_0_oe),
	.addq_0 /* IN */ (addq_0_[15:0]),
	.addq_1 /* IN */ (addq_1_[15:0]),
	.addq_2 /* IN */ (addq_2_[15:0]),
	.addq_3 /* IN */ (addq_3_[15:0]),
	.big_pix /* IN */ (big_pix),
	.dstdlo /* IN */ (dstdlo_[31:0]),
	.dstdhi /* IN */ (dstdhi_[31:0]),
	.dstzlo /* IN */ (dstzlo_[31:0]),
	.dstzhi /* IN */ (dstzhi_[31:0]),
	.data_sel /* IN */ (data_sel[1:0]),
	.data_ena /* IN */ (data_ena),
	.dstart /* IN */ (dstart[5:0]),
	.dend /* IN */ (dend[5:0]),
	.dbinh_n /* IN */ (dbinh_n[7:0]),
	.lfu_0 /* IN */ (lfu_0_[31:0]),
	.lfu_1 /* IN */ (lfu_1_[31:0]),
	.patd_0 /* IN */ (patd_0_[31:0]),
	.patd_1 /* IN */ (patd_1_[31:0]),
	.phrase_mode /* IN */ (phrase_mode),
	.srczlo /* IN */ (srczlo_[31:0]),
	.srczhi /* IN */ (srczhi_[31:0])
);
endmodule
