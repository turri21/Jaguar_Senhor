/* verilator lint_off LITENDIAN */
//`include "defs.v"

module j_fa23
(
	output s_0,
	output s_1,
	output s_2,
	output s_3,
	output s_4,
	output s_5,
	output s_6,
	output s_7,
	output s_8,
	output s_9,
	output s_10,
	output s_11,
	output s_12,
	output s_13,
	output s_14,
	output s_15,
	output s_16,
	output s_17,
	output s_18,
	output s_19,
	output s_20,
	output s_21,
	output s_22,
	input a_0,
	input a_1,
	input a_2,
	input a_3,
	input a_4,
	input a_5,
	input a_6,
	input a_7,
	input a_8,
	input a_9,
	input a_10,
	input a_11,
	input a_12,
	input a_13,
	input a_14,
	input a_15,
	input a_16,
	input a_17,
	input a_18,
	input a_19,
	input a_20,
	input a_21,
	input a_22,
	input b_0,
	input b_1,
	input b_2,
	input b_3,
	input b_4,
	input b_5,
	input b_6,
	input b_7,
	input b_8,
	input b_9,
	input b_10,
	input b_11,
	input b_12,
	input b_13,
	input b_14,
	input b_15,
	input b_16,
	input b_17,
	input b_18,
	input b_19,
	input b_20,
	input b_21,
	input b_22
);
wire zero;
wire s_23;
wire s_24;
wire s_25;
wire s_26;
wire s_27;
wire s_28;
wire s_29;
wire s_30;
wire s_31;
wire unused_0;
wire unused_1;
wire unused_2;

// DSP_F-35.NET (362) - zero : tie0
assign zero = 1'b0;

// DSP_F-35.NET (363) - fa32 : fa32
fa32 fa32_inst
(
	.s0 /* OUT */ (s_0),
	.s1 /* OUT */ (s_1),
	.s2 /* OUT */ (s_2),
	.s3 /* OUT */ (s_3),
	.s4 /* OUT */ (s_4),
	.s5 /* OUT */ (s_5),
	.s6 /* OUT */ (s_6),
	.s7 /* OUT */ (s_7),
	.s8 /* OUT */ (s_8),
	.s9 /* OUT */ (s_9),
	.s10 /* OUT */ (s_10),
	.s11 /* OUT */ (s_11),
	.s12 /* OUT */ (s_12),
	.s13 /* OUT */ (s_13),
	.s14 /* OUT */ (s_14),
	.s15 /* OUT */ (s_15),
	.s16 /* OUT */ (s_16),
	.s17 /* OUT */ (s_17),
	.s18 /* OUT */ (s_18),
	.s19 /* OUT */ (s_19),
	.s20 /* OUT */ (s_20),
	.s21 /* OUT */ (s_21),
	.s22 /* OUT */ (s_22),
	.s23 /* OUT */ (s_23),
	.s24 /* OUT */ (s_24),
	.s25 /* OUT */ (s_25),
	.s26 /* OUT */ (s_26),
	.s27 /* OUT */ (s_27),
	.s28 /* OUT */ (s_28),
	.s29 /* OUT */ (s_29),
	.s30 /* OUT */ (s_30),
	.s31 /* OUT */ (s_31),
	.co32 /* OUT */ (unused_0),
	.co31 /* OUT */ (unused_1),
	.co24 /* OUT */ (unused_2),
	.ci /* IN */ (zero),
	.a0 /* IN */ (a_0),
	.b0 /* IN */ (b_0),
	.a1 /* IN */ (a_1),
	.b1 /* IN */ (b_1),
	.a2 /* IN */ (a_2),
	.b2 /* IN */ (b_2),
	.a3 /* IN */ (a_3),
	.b3 /* IN */ (b_3),
	.a4 /* IN */ (a_4),
	.b4 /* IN */ (b_4),
	.a5 /* IN */ (a_5),
	.b5 /* IN */ (b_5),
	.a6 /* IN */ (a_6),
	.b6 /* IN */ (b_6),
	.a7 /* IN */ (a_7),
	.b7 /* IN */ (b_7),
	.a8 /* IN */ (a_8),
	.b8 /* IN */ (b_8),
	.a9 /* IN */ (a_9),
	.b9 /* IN */ (b_9),
	.a10 /* IN */ (a_10),
	.b10 /* IN */ (b_10),
	.a11 /* IN */ (a_11),
	.b11 /* IN */ (b_11),
	.a12 /* IN */ (a_12),
	.b12 /* IN */ (b_12),
	.a13 /* IN */ (a_13),
	.b13 /* IN */ (b_13),
	.a14 /* IN */ (a_14),
	.b14 /* IN */ (b_14),
	.a15 /* IN */ (a_15),
	.b15 /* IN */ (b_15),
	.a16 /* IN */ (a_16),
	.b16 /* IN */ (b_16),
	.a17 /* IN */ (a_17),
	.b17 /* IN */ (b_17),
	.a18 /* IN */ (a_18),
	.b18 /* IN */ (b_18),
	.a19 /* IN */ (a_19),
	.b19 /* IN */ (b_19),
	.a20 /* IN */ (a_20),
	.b20 /* IN */ (b_20),
	.a21 /* IN */ (a_21),
	.b21 /* IN */ (b_21),
	.a22 /* IN */ (a_22),
	.b22 /* IN */ (b_22),
	.a23 /* IN */ (zero),
	.b23 /* IN */ (zero),
	.a24 /* IN */ (zero),
	.b24 /* IN */ (zero),
	.a25 /* IN */ (zero),
	.b25 /* IN */ (zero),
	.a26 /* IN */ (zero),
	.b26 /* IN */ (zero),
	.a27 /* IN */ (zero),
	.b27 /* IN */ (zero),
	.a28 /* IN */ (zero),
	.b28 /* IN */ (zero),
	.a29 /* IN */ (zero),
	.b29 /* IN */ (zero),
	.a30 /* IN */ (zero),
	.b30 /* IN */ (zero),
	.a31 /* IN */ (zero),
	.b31 /* IN */ (zero)
);

// DSP_F-35.NET (372) - dummy[0-2] : dummy

// DSP_F-35.NET (373) - dummy[23-31] : dummy
endmodule
/* verilator lint_on LITENDIAN */
