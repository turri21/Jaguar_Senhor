//`include "defs.v"
// altera message_off 10036

module mem
(
	input bbreq_0,
	input bbreq_1,
	input gbreq_0,
	input gbreq_1,
	input obbreq,
	input sizin_0,
	input sizin_1,
	input dbrl_0,
	input dbrl_1,
	input dreqin,
	input rwin,
	input bs_0,
	input bs_1,
	input bs_2,
	input bs_3,
	input match,
	input intdev,
	input dram,
	input fextdev,
	input fintdev,
	input fdram,
	input from,
	input cpu32,
	input refreq,
	input dspd_0,
	input dspd_1,
	input romspd_0,
	input romspd_1,
	input iospd_0,
	input iospd_1,
	input a_0,
	input a_1,
	input a_2,
	input mw_0,
	input mw_1,
	input ourack,
	input resetl,
	input clk,
	input vcc,
	input gnd,
	input bglin,
	input brlin,
	input ihandler,
	input bigend,
	input bgain,
	input abs_2,
	input abs_3,
	input testen,
	input waitl,
	input fastrom,
	input m68k,
	input pclk,
	output ack,
	output bback,
	output gback,
	output obback,
	output romcsl_0,
	output romcsl_1,
	output rasl_0,
	output rasl_1,
	output casl_0,
	output casl_1,
	output oel_0,
	output oel_1,
	output oel_2,
	output wel_0,
	output wel_1,
	output wel_2,
	output wel_3,
	output wel_4,
	output wel_5,
	output wel_6,
	output wel_7,
	output sizout_0,
	output sizout_1,
	output sizout_2,
	output den_0,
	output den_1,
	output den_2,
	output aen,
	output dtackl,
	output brlout,
	output dbgl,
	output dreqlout,
	output d7a,
	output readt,
	output dinlatch_0,
	output dinlatch_1,
	output dinlatch_2,
	output dinlatch_3,
	output dinlatch_4,
	output dinlatch_5,
	output dinlatch_6,
	output dinlatch_7,
	output dmuxu_0,
	output dmuxu_1,
	output dmuxu_2,
	output dmuxd_0,
	output dmuxd_1,
	output dmuxd_2,
	output dren,
	output xdsrc,
	output maska_0,
	output maska_1,
	output maska_2,
	output at_0,
	output at_1,
	output at_2,
	output ainen,
	output newrow,
	output resrow,
	output mux,
	output refack,
	output reads,
	output wet,
	output oet,
	output ba,
	output intswe,
	output intwe,
	output dspcsl,
	output w_0_out,
	output w_0_oe,
	input w_0_in,
	output w_1_out,
	output w_1_oe,
	input w_1_in,
	output w_2_out,
	output w_2_oe,
	input w_2_in,
	output w_3_out,
	output w_3_oe,
	input w_3_in,
	output rw_out,
	output rw_oe,
	input rw_in,
	output mreq_out,
	output mreq_oe,
	input mreq_in,
	output justify_out,
	output justify_oe,
	input justify_in,
	input tlw,
	input ram_rdy,
	input sys_clk, // Generated
	
	output startcas_out
);
wire [1:0] bbreq = {bbreq_1,bbreq_0};
wire [1:0] gbreq = {gbreq_1,gbreq_0};
wire [1:0] sizin = {sizin_1,sizin_0};
wire [1:0] dbrl = {dbrl_1,dbrl_0};
wire [3:0] bs = {bs_3,bs_2,bs_1,bs_0};
wire [1:0] dspd = {dspd_1,dspd_0};
wire [1:0] romspd = {romspd_1,romspd_0};
wire [1:0] iospd = {iospd_1,iospd_0};
wire [2:0] a = {a_2,a_1,a_0};
wire [1:0] mw = {mw_1,mw_0};
wire [3:2] abs = {abs_3,abs_2};
wire [1:0] romcsl;
assign {romcsl_1,romcsl_0} = romcsl[1:0];
wire [1:0] rasl;
assign {rasl_1,rasl_0} = rasl[1:0];
wire [1:0] casl;
assign {casl_1,casl_0} = casl[1:0];
wire [2:0] oel;
assign {oel_2,oel_1,oel_0} = oel[2:0];
wire [7:0] wel;
assign {wel_7,wel_6,wel_5,wel_4,wel_3,wel_2,wel_1,wel_0} = wel[7:0];
wire [2:0] sizout;
assign {sizout_2,sizout_1,sizout_0} = sizout[2:0];
wire [2:0] den;
assign {den_2,den_1,den_0} = den[2:0];
wire [7:0] dinlatch;
assign {dinlatch_7,dinlatch_6,dinlatch_5,dinlatch_4,dinlatch_3,dinlatch_2,dinlatch_1,dinlatch_0} = dinlatch[7:0];
wire [2:0] dmuxu;
assign {dmuxu_2,dmuxu_1,dmuxu_0} = dmuxu[2:0];
wire [2:0] dmuxd;
assign {dmuxd_2,dmuxd_1,dmuxd_0} = dmuxd[2:0];
wire [2:0] maska;
assign {maska_2,maska_1,maska_0} = maska[2:0];
wire [2:0] at;
assign {at_2,at_1,at_0} = at[2:0];
wire [3:0] w_out;
assign {w_3_out,w_2_out,w_1_out,w_0_out} = w_out[3:0];
assign {w_3_oe,w_2_oe,w_1_oe} = {3{w_0_oe}};
wire [3:0] w_in = {w_3_in,w_2_in,w_1_in,w_0_in};
_mem mem_inst
(
	.bbreq /* IN */ (bbreq[1:0]),
	.gbreq /* IN */ (gbreq[1:0]),
	.obbreq /* IN */ (obbreq),
	.sizin /* IN */ (sizin[1:0]),
	.dbrl /* IN */ (dbrl[1:0]),
	.dreqin /* IN */ (dreqin),
	.rwin /* IN */ (rwin),
	.bs /* IN */ (bs[3:0]),
	.match /* IN */ (match),
	.intdev /* IN */ (intdev),
	.dram /* IN */ (dram),
	.fextdev /* IN */ (fextdev),
	.fintdev /* IN */ (fintdev),
	.fdram /* IN */ (fdram),
	.from /* IN */ (from),
	.cpu32 /* IN */ (cpu32),
	.refreq /* IN */ (refreq),
	.dspd /* IN */ (dspd[1:0]),
	.romspd /* IN */ (romspd[1:0]),
	.iospd /* IN */ (iospd[1:0]),
	.a /* IN */ (a[2:0]),
	.mw /* IN */ (mw[1:0]),
	.ourack /* IN */ (ourack),
	.resetl /* IN */ (resetl),
	.clk /* IN */ (clk),
	.bglin /* IN */ (bglin),
	.brlin /* IN */ (brlin),
	.ihandler /* IN */ (ihandler),
	.bigend /* IN */ (bigend),
	.bgain /* IN */ (bgain),
	.abs /* IN */ (abs[3:2]),
	.testen /* IN */ (testen),
	.waitl /* IN */ (waitl),
	.fastrom /* IN */ (fastrom),
	.m68k /* IN */ (m68k),
	.pclk /* IN */ (pclk),
	.ack /* OUT */ (ack),
	.bback /* OUT */ (bback),
	.gback /* OUT */ (gback),
	.obback /* OUT */ (obback),
	.romcsl /* OUT */ (romcsl[1:0]),
	.rasl /* OUT */ (rasl[1:0]),
	.casl /* OUT */ (casl[1:0]),
	.oel /* OUT */ (oel[2:0]),
	.wel /* OUT */ (wel[7:0]),
	.sizout /* OUT */ (sizout[2:0]),
	.den /* OUT */ (den[2:0]),
	.aen /* OUT */ (aen),
	.dtackl /* OUT */ (dtackl),
	.brlout /* OUT */ (brlout),
	.dbgl /* OUT */ (dbgl),
	.dreqlout /* OUT */ (dreqlout),
	.d7a /* OUT */ (d7a),
	.readt /* OUT */ (readt),
	.dinlatch /* OUT */ (dinlatch[7:0]),
	.dmuxu /* OUT */ (dmuxu[2:0]),
	.dmuxd /* OUT */ (dmuxd[2:0]),
	.dren /* OUT */ (dren),
	.xdsrc /* OUT */ (xdsrc),
	.maska /* OUT */ (maska[2:0]),
	.at /* OUT */ (at[2:0]),
	.ainen /* OUT */ (ainen),
	.newrow /* OUT */ (newrow),
	.resrow /* OUT */ (resrow),
	.mux /* OUT */ (mux),
	.refack /* OUT */ (refack),
	.reads /* OUT */ (reads),
	.wet /* OUT */ (wet),
	.oet /* OUT */ (oet),
	.ba /* OUT */ (ba),
	.intswe /* OUT */ (intswe),
	.intwe /* OUT */ (intwe),
	.dspcsl /* OUT */ (dspcsl),
	.w_out /* BUS */ (w_out[3:0]),
	.w_oe /* BUS */ (w_0_oe),
	.w_in /* BUS */ (w_in[3:0]),
	.rw_out /* BUS */ (rw_out),
	.rw_oe /* BUS */ (rw_oe),
	.rw_in /* BUS */ (rw_in),
	.mreq_out /* BUS */ (mreq_out),
	.mreq_oe /* BUS */ (mreq_oe),
	.mreq_in /* BUS */ (mreq_in),
	.justify_out /* BUS */ (justify_out),
	.justify_oe /* BUS */ (justify_oe),
	.justify_in /* BUS */ (justify_in),
	.tlw /* IN */ (tlw),
	.ram_rdy /* IN */ (ram_rdy),
	.sys_clk(sys_clk), // Generated
	.startcas_out(startcas_out)
);
endmodule
