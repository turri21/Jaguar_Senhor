//`include "defs.v"
// altera message_off 10036

module dbus
(
	input din_0,
	input din_1,
	input din_2,
	input din_3,
	input din_4,
	input din_5,
	input din_6,
	input din_7,
	input din_8,
	input din_9,
	input din_10,
	input din_11,
	input din_12,
	input din_13,
	input din_14,
	input din_15,
	input din_16,
	input din_17,
	input din_18,
	input din_19,
	input din_20,
	input din_21,
	input din_22,
	input din_23,
	input din_24,
	input din_25,
	input din_26,
	input din_27,
	input din_28,
	input din_29,
	input din_30,
	input din_31,
	input din_32,
	input din_33,
	input din_34,
	input din_35,
	input din_36,
	input din_37,
	input din_38,
	input din_39,
	input din_40,
	input din_41,
	input din_42,
	input din_43,
	input din_44,
	input din_45,
	input din_46,
	input din_47,
	input din_48,
	input din_49,
	input din_50,
	input din_51,
	input din_52,
	input din_53,
	input din_54,
	input din_55,
	input din_56,
	input din_57,
	input din_58,
	input din_59,
	input din_60,
	input din_61,
	input din_62,
	input din_63,
	input dr_0,
	input dr_1,
	input dr_2,
	input dr_3,
	input dr_4,
	input dr_5,
	input dr_6,
	input dr_7,
	input dr_8,
	input dr_9,
	input dr_10,
	input dr_11,
	input dr_12,
	input dr_13,
	input dr_14,
	input dr_15,
	input dinlatch_0,
	input dinlatch_1,
	input dinlatch_2,
	input dinlatch_3,
	input dinlatch_4,
	input dinlatch_5,
	input dinlatch_6,
	input dinlatch_7,
	input dmuxd_0,
	input dmuxd_1,
	input dmuxd_2,
	input dmuxu_0,
	input dmuxu_1,
	input dmuxu_2,
	input dren,
	input xdsrc,
	input ourack,
	input wd_0,
	input wd_1,
	input wd_2,
	input wd_3,
	input wd_4,
	input wd_5,
	input wd_6,
	input wd_7,
	input wd_8,
	input wd_9,
	input wd_10,
	input wd_11,
	input wd_12,
	input wd_13,
	input wd_14,
	input wd_15,
	input wd_16,
	input wd_17,
	input wd_18,
	input wd_19,
	input wd_20,
	input wd_21,
	input wd_22,
	input wd_23,
	input wd_24,
	input wd_25,
	input wd_26,
	input wd_27,
	input wd_28,
	input wd_29,
	input wd_30,
	input wd_31,
	input wd_32,
	input wd_33,
	input wd_34,
	input wd_35,
	input wd_36,
	input wd_37,
	input wd_38,
	input wd_39,
	input wd_40,
	input wd_41,
	input wd_42,
	input wd_43,
	input wd_44,
	input wd_45,
	input wd_46,
	input wd_47,
	input wd_48,
	input wd_49,
	input wd_50,
	input wd_51,
	input wd_52,
	input wd_53,
	input wd_54,
	input wd_55,
	input wd_56,
	input wd_57,
	input wd_58,
	input wd_59,
	input wd_60,
	input wd_61,
	input wd_62,
	input wd_63,
	input clk,
	output dp_0,
	output dp_1,
	output dp_2,
	output dp_3,
	output dp_4,
	output dp_5,
	output dp_6,
	output dp_7,
	output dp_8,
	output dp_9,
	output dp_10,
	output dp_11,
	output dp_12,
	output dp_13,
	output dp_14,
	output dp_15,
	output dob_0,
	output dob_1,
	output dob_2,
	output dob_3,
	output dob_4,
	output dob_5,
	output dob_6,
	output dob_7,
	output dob_8,
	output dob_9,
	output dob_10,
	output dob_11,
	output dob_12,
	output dob_13,
	output dob_14,
	output dob_15,
	output dout_16,
	output dout_17,
	output dout_18,
	output dout_19,
	output dout_20,
	output dout_21,
	output dout_22,
	output dout_23,
	output dout_24,
	output dout_25,
	output dout_26,
	output dout_27,
	output dout_28,
	output dout_29,
	output dout_30,
	output dout_31,
	output d5_32,
	output d5_33,
	output d5_34,
	output d5_35,
	output d5_36,
	output d5_37,
	output d5_38,
	output d5_39,
	output d5_40,
	output d5_41,
	output d5_42,
	output d5_43,
	output d5_44,
	output d5_45,
	output d5_46,
	output d5_47,
	output d5_48,
	output d5_49,
	output d5_50,
	output d5_51,
	output d5_52,
	output d5_53,
	output d5_54,
	output d5_55,
	output d5_56,
	output d5_57,
	output d5_58,
	output d5_59,
	output d5_60,
	output d5_61,
	output d5_62,
	output d5_63,
	output d_0,
	output d_1,
	output d_2,
	output d_3,
	output d_4,
	output d_5,
	output d_6,
	output d_7,
	output d_8,
	output d_9,
	output d_10,
	output d_11,
	output d_12,
	output d_13,
	output d_14,
	output d_15,
	output d_16,
	output d_17,
	output d_18,
	output d_19,
	output d_20,
	output d_21,
	output d_22,
	output d_23,
	output d_24,
	output d_25,
	output d_26,
	output d_27,
	output d_28,
	output d_29,
	output d_30,
	output d_31,
	output d_32,
	output d_33,
	output d_34,
	output d_35,
	output d_36,
	output d_37,
	output d_38,
	output d_39,
	output d_40,
	output d_41,
	output d_42,
	output d_43,
	output d_44,
	output d_45,
	output d_46,
	output d_47,
	output d_48,
	output d_49,
	output d_50,
	output d_51,
	output d_52,
	output d_53,
	output d_54,
	output d_55,
	output d_56,
	output d_57,
	output d_58,
	output d_59,
	output d_60,
	output d_61,
	output d_62,
	output d_63,
	input sys_clk // Generated
);

wire [63:0] din = {din_63,din_62,din_61,din_60,
din_59,din_58,din_57,din_56,din_55,din_54,din_53,din_52,din_51,din_50,
din_49,din_48,din_47,din_46,din_45,din_44,din_43,din_42,din_41,din_40,
din_39,din_38,din_37,din_36,din_35,din_34,din_33,din_32,din_31,din_30,
din_29,din_28,din_27,din_26,din_25,din_24,din_23,din_22,din_21,din_20,
din_19,din_18,din_17,din_16,din_15,din_14,din_13,din_12,din_11,din_10,
din_9,din_8,din_7,din_6,din_5,din_4,din_3,din_2,din_1,din_0};
wire [15:0] dr = {dr_15,dr_14,dr_13,dr_12,dr_11,dr_10,
dr_9,dr_8,dr_7,dr_6,dr_5,dr_4,dr_3,dr_2,dr_1,dr_0};
wire [7:0] dinlatch = {dinlatch_7,dinlatch_6,dinlatch_5,dinlatch_4,dinlatch_3,dinlatch_2,dinlatch_1,dinlatch_0};
wire [2:0] dmuxd = {dmuxd_2,dmuxd_1,dmuxd_0};
wire [2:0] dmuxu = {dmuxu_2,dmuxu_1,dmuxu_0};
wire [63:0] wd = {wd_63,wd_62,wd_61,wd_60,
wd_59,wd_58,wd_57,wd_56,wd_55,wd_54,wd_53,wd_52,wd_51,wd_50,
wd_49,wd_48,wd_47,wd_46,wd_45,wd_44,wd_43,wd_42,wd_41,wd_40,
wd_39,wd_38,wd_37,wd_36,wd_35,wd_34,wd_33,wd_32,wd_31,wd_30,
wd_29,wd_28,wd_27,wd_26,wd_25,wd_24,wd_23,wd_22,wd_21,wd_20,
wd_19,wd_18,wd_17,wd_16,wd_15,wd_14,wd_13,wd_12,wd_11,wd_10,
wd_9,wd_8,wd_7,wd_6,wd_5,wd_4,wd_3,wd_2,wd_1,wd_0};
wire [15:0] dp;
assign {dp_15,dp_14,dp_13,dp_12,dp_11,dp_10,
dp_9,dp_8,dp_7,dp_6,dp_5,dp_4,dp_3,dp_2,dp_1,dp_0} = dp[15:0];
wire [15:0] dob;
assign {dob_15,dob_14,dob_13,dob_12,dob_11,dob_10,
dob_9,dob_8,dob_7,dob_6,dob_5,dob_4,dob_3,dob_2,dob_1,dob_0} = dob[15:0];
wire [31:16] dout;
assign {dout_31,dout_30,
dout_29,dout_28,dout_27,dout_26,dout_25,dout_24,dout_23,dout_22,dout_21,dout_20,
dout_19,dout_18,dout_17,dout_16} = dout[31:16];
wire [63:32] d5;
assign {d5_63,d5_62,d5_61,d5_60,
d5_59,d5_58,d5_57,d5_56,d5_55,d5_54,d5_53,d5_52,d5_51,d5_50,
d5_49,d5_48,d5_47,d5_46,d5_45,d5_44,d5_43,d5_42,d5_41,d5_40,
d5_39,d5_38,d5_37,d5_36,d5_35,d5_34,d5_33,d5_32} = d5[63:32];
wire [63:0] d;
assign {d_63,d_62,d_61,d_60,
d_59,d_58,d_57,d_56,d_55,d_54,d_53,d_52,d_51,d_50,
d_49,d_48,d_47,d_46,d_45,d_44,d_43,d_42,d_41,d_40,
d_39,d_38,d_37,d_36,d_35,d_34,d_33,d_32,d_31,d_30,
d_29,d_28,d_27,d_26,d_25,d_24,d_23,d_22,d_21,d_20,
d_19,d_18,d_17,d_16,d_15,d_14,d_13,d_12,d_11,d_10,
d_9,d_8,d_7,d_6,d_5,d_4,d_3,d_2,d_1,d_0} = d[63:0];
// TOM.NET (363) - dbus : dbus
_dbus dbus_inst
(
	.din /* IN */ (din[63:0]),
	.dr /* IN */ (dr[15:0]),
	.dinlatch /* IN */ (dinlatch[7:0]),
	.dmuxd /* IN */ (dmuxd[2:0]),
	.dmuxu /* IN */ (dmuxu[2:0]),
	.dren /* IN */ (dren),
	.xdsrc /* IN */ (xdsrc),
	.ourack /* IN */ (ourack),
	.wd /* IN */ (wd[63:0]),
	.clk /* IN */ (clk),
	.dp /* OUT */ (dp[15:0]),
	.dob /* OUT */ (dob[15:0]),
	.dout /* OUT */ (dout[31:16]),
	.d5 /* OUT */ (d5[63:32]),
	.d /* OUT */ (d[63:0]),
	.sys_clk(sys_clk) // Generated
);
endmodule
