module j_jerry
(
	input xdspcsl,
	input xpclkosc,
	input xpclkin,
	input xdbgl,
	input xoel_0,
	input xwel_0,
	input xserin,
	input xdtackl,
	input xi2srxd,
	input xeint_0,
	input xeint_1,
	input xtest,
	input xchrin,
	input xresetil,
	output xd_0_out,
	output xd_0_oe,
	input xd_0_in,
	output xd_1_out,
	output xd_1_oe,
	input xd_1_in,
	output xd_2_out,
	output xd_2_oe,
	input xd_2_in,
	output xd_3_out,
	output xd_3_oe,
	input xd_3_in,
	output xd_4_out,
	output xd_4_oe,
	input xd_4_in,
	output xd_5_out,
	output xd_5_oe,
	input xd_5_in,
	output xd_6_out,
	output xd_6_oe,
	input xd_6_in,
	output xd_7_out,
	output xd_7_oe,
	input xd_7_in,
	output xd_8_out,
	output xd_8_oe,
	input xd_8_in,
	output xd_9_out,
	output xd_9_oe,
	input xd_9_in,
	output xd_10_out,
	output xd_10_oe,
	input xd_10_in,
	output xd_11_out,
	output xd_11_oe,
	input xd_11_in,
	output xd_12_out,
	output xd_12_oe,
	input xd_12_in,
	output xd_13_out,
	output xd_13_oe,
	input xd_13_in,
	output xd_14_out,
	output xd_14_oe,
	input xd_14_in,
	output xd_15_out,
	output xd_15_oe,
	input xd_15_in,
	output xd_16_out,
	output xd_16_oe,
	input xd_16_in,
	output xd_17_out,
	output xd_17_oe,
	input xd_17_in,
	output xd_18_out,
	output xd_18_oe,
	input xd_18_in,
	output xd_19_out,
	output xd_19_oe,
	input xd_19_in,
	output xd_20_out,
	output xd_20_oe,
	input xd_20_in,
	output xd_21_out,
	output xd_21_oe,
	input xd_21_in,
	output xd_22_out,
	output xd_22_oe,
	input xd_22_in,
	output xd_23_out,
	output xd_23_oe,
	input xd_23_in,
	output xd_24_out,
	output xd_24_oe,
	input xd_24_in,
	output xd_25_out,
	output xd_25_oe,
	input xd_25_in,
	output xd_26_out,
	output xd_26_oe,
	input xd_26_in,
	output xd_27_out,
	output xd_27_oe,
	input xd_27_in,
	output xd_28_out,
	output xd_28_oe,
	input xd_28_in,
	output xd_29_out,
	output xd_29_oe,
	input xd_29_in,
	output xd_30_out,
	output xd_30_oe,
	input xd_30_in,
	output xd_31_out,
	output xd_31_oe,
	input xd_31_in,
	output xa_0_out,
	output xa_0_oe,
	input xa_0_in,
	output xa_1_out,
	output xa_1_oe,
	input xa_1_in,
	output xa_2_out,
	output xa_2_oe,
	input xa_2_in,
	output xa_3_out,
	output xa_3_oe,
	input xa_3_in,
	output xa_4_out,
	output xa_4_oe,
	input xa_4_in,
	output xa_5_out,
	output xa_5_oe,
	input xa_5_in,
	output xa_6_out,
	output xa_6_oe,
	input xa_6_in,
	output xa_7_out,
	output xa_7_oe,
	input xa_7_in,
	output xa_8_out,
	output xa_8_oe,
	input xa_8_in,
	output xa_9_out,
	output xa_9_oe,
	input xa_9_in,
	output xa_10_out,
	output xa_10_oe,
	input xa_10_in,
	output xa_11_out,
	output xa_11_oe,
	input xa_11_in,
	output xa_12_out,
	output xa_12_oe,
	input xa_12_in,
	output xa_13_out,
	output xa_13_oe,
	input xa_13_in,
	output xa_14_out,
	output xa_14_oe,
	input xa_14_in,
	output xa_15_out,
	output xa_15_oe,
	input xa_15_in,
	output xa_16_out,
	output xa_16_oe,
	input xa_16_in,
	output xa_17_out,
	output xa_17_oe,
	input xa_17_in,
	output xa_18_out,
	output xa_18_oe,
	input xa_18_in,
	output xa_19_out,
	output xa_19_oe,
	input xa_19_in,
	output xa_20_out,
	output xa_20_oe,
	input xa_20_in,
	output xa_21_out,
	output xa_21_oe,
	input xa_21_in,
	output xa_22_out,
	output xa_22_oe,
	input xa_22_in,
	output xa_23_out,
	output xa_23_oe,
	input xa_23_in,
	output xjoy_0_out,
	output xjoy_0_oe,
	input xjoy_0_in,
	output xjoy_1_out,
	output xjoy_1_oe,
	input xjoy_1_in,
	output xjoy_2_out,
	output xjoy_2_oe,
	input xjoy_2_in,
	output xjoy_3_out,
	output xjoy_3_oe,
	input xjoy_3_in,
	output xgpiol_0_out,
	output xgpiol_0_oe,
	input xgpiol_0_in,
	output xgpiol_1_out,
	output xgpiol_1_oe,
	input xgpiol_1_in,
	output xgpiol_2_out,
	output xgpiol_2_oe,
	input xgpiol_2_in,
	output xgpiol_3_out,
	output xgpiol_3_oe,
	input xgpiol_3_in,
	output xsck_out,
	output xsck_oe,
	input xsck_in,
	output xws_out,
	output xws_oe,
	input xws_in,
	output xvclk_out,
	output xvclk_oe,
	input xvclk_in,
	output xsiz_0_out,
	output xsiz_0_oe,
	input xsiz_0_in,
	output xsiz_1_out,
	output xsiz_1_oe,
	input xsiz_1_in,
	output xrw_out,
	output xrw_oe,
	input xrw_in,
	output xdreql_out,
	output xdreql_oe,
	input xdreql_in,
	output xdbrl_0,
	output xdbrl_1,
	output xint,
	output xserout,
	output xgpiol_4,
	output xgpiol_5,
	output xvclkdiv,
	output xchrdiv,
	output xpclkout,
	output xpclkdiv,
	output xresetl,
	output xchrout,
	output xrdac_0,
	output xrdac_1,
	output xldac_0,
	output xldac_1,
	output xiordl,
	output xiowrl,
	output xi2stxd,
	output xcpuclk,
	input tlw,
	input tlw_0,
	input tlw_1,
	input tlw_2,
	output aen,
	output den,
	output ainen,
	output [15:0] snd_l,
	output [15:0] snd_r,
	output snd_l_en,
	output snd_r_en,
	output snd_clk,
	
	output [15:0] dspwd,
	
	input sys_clk // Generated
);
wire [1:0] xeint = {xeint_1,xeint_0};
wire [31:0] xd_out; //
assign {xd_31_out,xd_30_out,
xd_29_out,xd_28_out,xd_27_out,xd_26_out,xd_25_out,xd_24_out,xd_23_out,xd_22_out,xd_21_out,xd_20_out,
xd_19_out,xd_18_out,xd_17_out,xd_16_out,xd_15_out,xd_14_out,xd_13_out,xd_12_out,xd_11_out,xd_10_out,
xd_9_out,xd_8_out,xd_7_out,xd_6_out,xd_5_out,xd_4_out,xd_3_out,xd_2_out,xd_1_out,xd_0_out} = xd_out[31:0];
wire [31:0] xd_oe;
assign {xd_31_oe,xd_30_oe,
xd_29_oe,xd_28_oe,xd_27_oe,xd_26_oe,xd_25_oe,xd_24_oe,xd_23_oe,xd_22_oe,xd_21_oe,xd_20_oe,
xd_19_oe,xd_18_oe,xd_17_oe,xd_16_oe,xd_15_oe,xd_14_oe,xd_13_oe,xd_12_oe,xd_11_oe,xd_10_oe,
xd_9_oe,xd_8_oe,xd_7_oe,xd_6_oe,xd_5_oe,xd_4_oe,xd_3_oe,xd_2_oe,xd_1_oe,xd_0_oe} = xd_oe[31:0];
wire [31:0] xd_in = {xd_31_in,xd_30_in,
xd_29_in,xd_28_in,xd_27_in,xd_26_in,xd_25_in,xd_24_in,xd_23_in,xd_22_in,xd_21_in,xd_20_in,
xd_19_in,xd_18_in,xd_17_in,xd_16_in,xd_15_in,xd_14_in,xd_13_in,xd_12_in,xd_11_in,xd_10_in,
xd_9_in,xd_8_in,xd_7_in,xd_6_in,xd_5_in,xd_4_in,xd_3_in,xd_2_in,xd_1_in,xd_0_in};
wire [23:0] xa_out; //
assign {xa_23_out,xa_22_out,xa_21_out,xa_20_out,
xa_19_out,xa_18_out,xa_17_out,xa_16_out,xa_15_out,xa_14_out,xa_13_out,xa_12_out,xa_11_out,xa_10_out,
xa_9_out,xa_8_out,xa_7_out,xa_6_out,xa_5_out,xa_4_out,xa_3_out,xa_2_out,xa_1_out,xa_0_out} = xa_out[23:0];
wire [23:0] xa_oe;
assign {xa_23_oe,xa_22_oe,xa_21_oe,xa_20_oe,
xa_19_oe,xa_18_oe,xa_17_oe,xa_16_oe,xa_15_oe,xa_14_oe,xa_13_oe,xa_12_oe,xa_11_oe,xa_10_oe,
xa_9_oe,xa_8_oe,xa_7_oe,xa_6_oe,xa_5_oe,xa_4_oe,xa_3_oe,xa_2_oe,xa_1_oe,xa_0_oe} = xa_oe[23:0];
wire [23:0] xa_in = {xa_23_in,xa_22_in,xa_21_in,xa_20_in,
xa_19_in,xa_18_in,xa_17_in,xa_16_in,xa_15_in,xa_14_in,xa_13_in,xa_12_in,xa_11_in,xa_10_in,
xa_9_in,xa_8_in,xa_7_in,xa_6_in,xa_5_in,xa_4_in,xa_3_in,xa_2_in,xa_1_in,xa_0_in};
wire [3:0] xjoy_out; //
assign {xjoy_3_out,xjoy_2_out,xjoy_1_out,xjoy_0_out} = xjoy_out[3:0];
wire [3:0] xjoy_oe;
assign {xjoy_3_oe,xjoy_2_oe,xjoy_1_oe,xjoy_0_oe} = xjoy_oe[3:0];
wire [3:0] xjoy_in = {xjoy_3_in,xjoy_2_in,xjoy_1_in,xjoy_0_in};
wire [5:0] xgpiol_out; // 4 and 5 included
assign {xgpiol_5,xgpiol_4,xgpiol_3_out,xgpiol_2_out,xgpiol_1_out,xgpiol_0_out} = xgpiol_out[5:0];
wire [3:0] xgpiol_oe;
assign {xgpiol_3_oe,xgpiol_2_oe,xgpiol_1_oe,xgpiol_0_oe} = xgpiol_oe[3:0];
wire [3:0] xgpiol_in = {xgpiol_3_in,xgpiol_2_in,xgpiol_1_in,xgpiol_0_in};
wire [1:0] xsiz_out; //
assign {xsiz_1_out,xsiz_0_out} = xsiz_out[1:0];
wire [1:0] xsiz_oe;
assign {xsiz_1_oe,xsiz_0_oe} = xsiz_oe[1:0];
wire [1:0] xsiz_in = {xsiz_1_in,xsiz_0_in};
wire [1:0] xdbrl; //
assign {xdbrl_1,xdbrl_0} = xdbrl[1:0];
wire [1:0] xrdac; //
assign {xrdac_1,xrdac_0} = xrdac[1:0];
wire [1:0] xldac; //
assign {xldac_1,xldac_0} = xldac[1:0];
_j_jerry jerry_inst
(
	.xdspcsl(xdspcsl),
	.xpclkosc(xpclkosc),
	.xpclkin(xpclkout),
	.xdbgl(xdbgl),
	.xoel_0(xoel_0),
	.xwel_0(xwel_0),
	.xserin(xserin),
	.xdtackl(xdtackl),
	.xi2srxd(xi2srxd),
	.xeint(xeint[1:0]),
	.xtest(xtest),
	.xchrin(xchrin), // Should be 14.3mhz, ntsc clock?
	.xresetil(xresetil),
	.xd_out(xd_out[31:0]),
	.xd_oe(xd_oe[31:0]),
	.xd_in(xd_in[31:0]),
	.xa_out(xa_out[23:0]),
	.xa_oe(xa_oe[23:0]),
	.xa_in(xa_in[23:0]),
	.xjoy_out(xjoy_out[3:0]),
	.xjoy_oe(xjoy_oe[3:0]),
	.xjoy_in(xjoy_in[3:0]),
	.xgpiol_out(xgpiol_out[5:0]),//4 and 5 included
	.xgpiol_oe(xgpiol_oe[3:0]),
	.xgpiol_in(xgpiol_in[3:0]),
	.xsck_out(xsck_out),
	.xsck_oe(xsck_oe),
	.xsck_in(xsck_in),
	.xws_out(xws_out),
	.xws_oe(xws_oe),
	.xws_in(xws_in),
	.xvclk_out(xvclk_out),
	.xvclk_oe(xvclk_oe),
	.xvclk_in(xvclk_in),
	.xsiz_out(xsiz_out[1:0]),
	.xsiz_oe(xsiz_oe[1:0]),
	.xsiz_in(xsiz_in[1:0]),
	.xrw_out(xrw_out),
	.xrw_oe(xrw_oe),
	.xrw_in(xrw_in),
	.xdreql_out(xdreql_out),
	.xdreql_oe(xdreql_oe),
	.xdreql_in(xdreql_in),
	.xdbrl(xdbrl[1:0]),
	.xint(xint),
	.xserout(xserout),
	.xvclkdiv(xvclkdiv),
	.xchrdiv(xchrdiv),
	.xpclkout(xpclkout),
	.xpclkdiv(xpclkdiv),
	.xresetl(xresetl),
	.xchrout(xchrout),
	.xrdac(xrdac[1:0]),
	.xldac(xldac[1:0]),
	.xiordl(xiordl),
	.xiowrl(xiowrl),
	.xi2stxd(xi2stxd),
	.xcpuclk(xcpuclk),
	.tlw(tlw),
	.tlw_0(tlw_0),
	.tlw_1(tlw_1),
	.tlw_2(tlw_2),
	//.tlw(xpclk), // /!\
	.aen(aen),
	.den(den),
	.ainen(ainen),
	.snd_l(snd_l[15:0]),
	.snd_r(snd_r[15:0]),
	.snd_l_en(snd_l_en),
	.snd_r_en(snd_r_en),
	.snd_clk(snd_clk),
	.dspwd( dspwd[15:0] ),

	.sys_clk(sys_clk)
);

endmodule
