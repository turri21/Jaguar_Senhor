module barrel32
(
	output z_0,
	output z_1,
	output z_2,
	output z_3,
	output z_4,
	output z_5,
	output z_6,
	output z_7,
	output z_8,
	output z_9,
	output z_10,
	output z_11,
	output z_12,
	output z_13,
	output z_14,
	output z_15,
	output z_16,
	output z_17,
	output z_18,
	output z_19,
	output z_20,
	output z_21,
	output z_22,
	output z_23,
	output z_24,
	output z_25,
	output z_26,
	output z_27,
	output z_28,
	output z_29,
	output z_30,
	output z_31,
	input mux_0,
	input mux_1,
	input sft_0,
	input sft_1,
	input sft_2,
	input sft_3,
	input sft_4,
	input flin,
	input a_0,
	input a_1,
	input a_2,
	input a_3,
	input a_4,
	input a_5,
	input a_6,
	input a_7,
	input a_8,
	input a_9,
	input a_10,
	input a_11,
	input a_12,
	input a_13,
	input a_14,
	input a_15,
	input a_16,
	input a_17,
	input a_18,
	input a_19,
	input a_20,
	input a_21,
	input a_22,
	input a_23,
	input a_24,
	input a_25,
	input a_26,
	input a_27,
	input a_28,
	input a_29,
	input a_30,
	input a_31
);
wire [31:0] z;
assign {z_31,z_30,
z_29,z_28,z_27,z_26,z_25,z_24,z_23,z_22,z_21,z_20,
z_19,z_18,z_17,z_16,z_15,z_14,z_13,z_12,z_11,z_10,
z_9,z_8,z_7,z_6,z_5,z_4,z_3,z_2,z_1,z_0} = z[31:0];
wire [1:0] mux = {mux_1,mux_0};
wire [4:0] sft = {sft_4,sft_3,sft_2,sft_1,sft_0};
wire [31:0] a = {a_31,a_30,
a_29,a_28,a_27,a_26,a_25,a_24,a_23,a_22,a_21,a_20,
a_19,a_18,a_17,a_16,a_15,a_14,a_13,a_12,a_11,a_10,
a_9,a_8,a_7,a_6,a_5,a_4,a_3,a_2,a_1,a_0};
_barrel32 brl_inst
(
	.z /* OUT */ (z[31:0]),
	.mux /* IN */ (mux[1:0]),
	.sft /* IN */ (sft[4:0]),
	.flin /* IN */ (flin),
	.a /* IN */ (a[31:0])
);
endmodule
